module	OR4(a, b, c, d, z);

input	a, b, c, d;
output	z;

or #1 g1(z, a, b, c, d);

endmodule
