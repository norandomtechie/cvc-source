module	AN5(a, b, c, d, e, z);

input	a, b, c, d, e;
output	z;

and #1 g1(z, a, b, c, d, e);

endmodule
