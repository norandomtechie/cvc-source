module 	BUF8A(a, z);

input   a;
output  z;

buf #1 g1(z, a);

endmodule
