// DA Solutions Ltd., Texas Instruments provided Multiplier benchmark
// Public domain Verilog coded gate level circuit
// Created 1-Sep-94, D. J. Wharton
// VHDL equivalent model also available
// Library used TI TGC1000_2.1 5v CMOS

module csa_mult_n17_m17_2

       ( A_16_port, A_15_port, A_14_port, A_13_port, A_12_port, A_11_port, 
         A_10_port, A_9_port, A_8_port, A_7_port, A_6_port, A_5_port, A_4_port,
         A_3_port, A_2_port, A_1_port, A_0_port, B_16_port, B_15_port, 
         B_14_port, B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, 
         B_8_port, B_7_port, B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, 
         B_1_port, B_0_port, CTL, PRODUCT_33_port, 
         PRODUCT_32_port, PRODUCT_31_port, PRODUCT_30_port, PRODUCT_29_port, 
         PRODUCT_28_port, PRODUCT_27_port, PRODUCT_26_port, PRODUCT_25_port, 
         PRODUCT_24_port, PRODUCT_23_port, PRODUCT_22_port, PRODUCT_21_port, 
         PRODUCT_20_port, PRODUCT_19_port, PRODUCT_18_port, PRODUCT_17_port, 
         PRODUCT_16_port, PRODUCT_15_port, PRODUCT_14_port, PRODUCT_13_port, 
         PRODUCT_12_port, PRODUCT_11_port, PRODUCT_10_port, PRODUCT_9_port, 
         PRODUCT_8_port, PRODUCT_7_port, PRODUCT_6_port, PRODUCT_5_port, 
         PRODUCT_4_port, PRODUCT_3_port, PRODUCT_2_port, PRODUCT_1_port, 
         PRODUCT_0_port );
   
input    A_16_port, A_15_port, A_14_port, A_13_port, A_12_port, A_11_port,
         A_10_port, A_9_port, A_8_port, A_7_port, A_6_port, A_5_port, A_4_port,
         A_3_port, A_2_port, A_1_port, A_0_port, B_16_port, B_15_port,
         B_14_port, B_13_port, B_12_port, B_11_port, B_10_port, B_9_port,
         B_8_port, B_7_port, B_6_port, B_5_port, B_4_port, B_3_port, B_2_port,
         B_1_port, B_0_port, CTL;

output   PRODUCT_33_port,
         PRODUCT_32_port, PRODUCT_31_port, PRODUCT_30_port, PRODUCT_29_port,
         PRODUCT_28_port, PRODUCT_27_port, PRODUCT_26_port, PRODUCT_25_port,
         PRODUCT_24_port, PRODUCT_23_port, PRODUCT_22_port, PRODUCT_21_port,
         PRODUCT_20_port, PRODUCT_19_port, PRODUCT_18_port, PRODUCT_17_port,
         PRODUCT_16_port, PRODUCT_15_port, PRODUCT_14_port, PRODUCT_13_port,
         PRODUCT_12_port, PRODUCT_11_port, PRODUCT_10_port, PRODUCT_9_port,
         PRODUCT_8_port, PRODUCT_7_port, PRODUCT_6_port, PRODUCT_5_port,
         PRODUCT_4_port, PRODUCT_3_port, PRODUCT_2_port, PRODUCT_1_port,
         PRODUCT_0_port;

wire  n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, 
      n4299, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, 
      n4379, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, 
      n4459, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, 
      n4539, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, 
      n4619, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, 
      n4189, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, 
      n4269, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, 
      n4349, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, 
      n4429, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, 
      n4509, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, 
      n4989, n5019, n5018, n5017, n5016, n5015, n5014, n5013, n5012, n5011, 
      n5010, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, 
      n4079, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, 
      n4159, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, 
      n4239, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, 
      n4319, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, 
      n4799, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, 
      n4879, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, 
      n4959, n5209, n5208, n5207, n5206, n5205, n5204, n5203, n5202, n5201, 
      n3980, n5200, n3981, n3982, n3983, n3984, n3985, n3986, n5129, n3987, 
      n5128, n3988, n5127, n3989, n5126, n5125, n5124, n5123, n5122, n5121, 
      n5120, n5049, n5048, n5047, n5046, n5045, n5044, n5043, n5042, n5041, 
      n5040, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, 
      n4049, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, 
      n4129, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, 
      n4209, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, 
      n4689, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, 
      n4769, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, 
      n4849, n4920, n4921, n4922, n4923, n3870, n4924, n3871, n4925, n3872, 
      n4926, n3873, n4927, n3874, n4928, n3875, n4929, n3876, n3877, n3878, 
      n3879, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n5159, n3957, 
      n5158, n3958, n5157, n3959, n5156, n5155, n5154, n5153, n5152, n5151, 
      n5150, n5079, n5078, n5077, n5076, n5075, n5074, n5073, n5072, n5071, 
      n5070, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
      n4019, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, 
      n4499, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, 
      n4579, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, 
      n4659, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, 
      n4739, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, 
      n4819, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n5189, n3927, 
      n5188, n3928, n5187, n3929, n5186, n5185, n5184, n5183, n5182, n5181, 
      n5180, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, 
      n4389, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, 
      n4469, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, 
      n4549, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, 
      n4629, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, 
      n4709, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, 
      n4199, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, 
      n4279, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, 
      n4359, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, 
      n4439, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, 
      n4519, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, 
      n4999, n5009, n5008, n5007, n5006, n5005, n5004, n5003, n5002, n5001, 
      n5000, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, 
      n4089, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, 
      n4169, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, 
      n4249, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, 
      n4329, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, 
      n4409, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, 
      n4889, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, 
      n4969, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n5119, n3997, 
      n5118, n3998, n5117, n3999, n5116, n5115, n5114, n5113, n5112, n5111, 
      n5110, n5039, n5038, n5037, n5036, n5035, n5034, n5033, n5032, n5031, 
      n5030, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, 
      n4059, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, 
      n4139, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, 
      n4219, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, 
      n4699, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, 
      n4779, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, 
      n4859, n4930, n4931, n4932, n4933, n3880, n4934, n3881, n4935, n3882, 
      n4936, n3883, n4937, n3884, n4938, n3885, n4939, n3886, n3887, n3888, 
      n3889, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n5149, n3967, 
      n5148, n3968, n5147, n3969, n5146, n5145, n5144, n5143, n5142, n5141, 
      n5140, n5069, n5068, n5067, n5066, n5065, n5064, n5063, n5062, n5061, 
      n5060, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, 
      n4029, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, 
      n4109, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, 
      n4589, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, 
      n4669, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, 
      n4749, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, 
      n4829, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, 
      n4909, n3858, n3859, n3930, n3931, n3932, n3933, n3934, n3935, n3936, 
      n5179, n3937, n5178, n3938, n5177, n3939, n5176, n5175, n5174, n5173, 
      n5172, n5171, n5170, n5099, n5098, n5097, n5096, n5095, n5094, n5093, 
      n5092, n5091, n5090, n4390, n4391, n4392, n4393, n4394, n4395, n4396, 
      n4397, n4398, n4399, n4470, n4471, n4472, n4473, n4474, n4475, n4476, 
      n4477, n4478, n4479, n4550, n4551, n4552, n4553, n4554, n4555, n4556, 
      n4557, n4558, n4559, n4630, n4631, n4632, n4633, n4634, n4635, n4636, 
      n4637, n4638, n4639, n4710, n4711, n4712, n4713, n4714, n4715, n4716, 
      n4717, n4718, n4719, n3900, n3901, n3902, n3903, n3904, n3905, n3906, 
      n3907, n3908, n3909, n4280, n4281, n4282, n4283, n4284, n4285, n4286, 
      n4287, n4288, n4289, n4360, n4361, n4362, n4363, n4364, n4365, n4366, 
      n4367, n4368, n4369, n4440, n4441, n4442, n4443, n4444, n4445, n4446, 
      n4447, n4448, n4449, n4520, n4521, n4522, n4523, n4524, n4525, n4526, 
      n4527, n4528, n4529, n4600, n4601, n4602, n4603, n4604, n4605, n4606, 
      n4607, n4608, n4609, n4090, n4091, n4092, n4093, n4094, n4095, n4096, 
      n4097, n4098, n4099, n4170, n4171, n4172, n4173, n4174, n4175, n4176, 
      n4177, n4178, n4179, n4250, n4251, n4252, n4253, n4254, n4255, n4256, 
      n4257, n4258, n4259, n4330, n4331, n4332, n4333, n4334, n4335, n4336, 
      n4337, n4338, n4339, n4410, n4411, n4412, n4413, n4414, n4415, n4416, 
      n4417, n4418, n4419, n4890, n4891, n4892, n4893, n4894, n4895, n4896, 
      n4897, n4898, n4899, n4970, n4971, n4972, n4973, n4974, n4975, n4976, 
      n4977, n4978, n4979, n5109, n5108, n5107, n5106, n5105, n5104, n5103, 
      n5102, n5101, n5100, n5029, n5028, n5027, n5026, n5025, n5024, n5023, 
      n5022, n5021, n5020, n4060, n4061, n4062, n4063, n4064, n4065, n4066, 
      n4067, n4068, n4069, n4140, n4141, n4142, n4143, n4144, n4145, n4146, 
      n4147, n4148, n4149, n4220, n4221, n4222, n4223, n4224, n4225, n4226, 
      n4227, n4228, n4229, n4300, n4301, n4302, n4303, n4304, n4305, n4306, 
      n4307, n4308, n4309, n4780, n4781, n4782, n4783, n4784, n4785, n4786, 
      n4787, n4788, n4789, n4860, n4861, n4862, n4863, n4864, n4865, n4866, 
      n4867, n4868, n4869, n4940, n4941, n4942, n4943, n3890, n4944, n3891, 
      n4945, n3892, n4946, n3893, n4947, n3894, n4948, n3895, n4949, n3896, 
      n3897, n5218, n3898, n5217, n3899, n5216, n5215, n5214, n5213, n5212, 
      n5211, n3970, n5210, n3971, n3972, n3973, n3974, n3975, n3976, n5139, 
      n3977, n5138, n3978, n5137, n3979, n5136, n5135, n5134, n5133, n5132, 
      n5131, n5130, n5059, n5058, n5057, n5056, n5055, n5054, n5053, n5052, 
      n5051, n5050, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, 
      n4038, n4039, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
      n4118, n4119, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, 
      n4598, n4599, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, 
      n4678, n4679, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, 
      n4758, n4759, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, 
      n4838, n4839, n4910, n4911, n4912, n4913, n3860, n4914, n3861, n4915, 
      n3862, n4916, n3863, n4917, n3864, n4918, n3865, n4919, n3866, n3867, 
      n3868, n3869, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n5169, 
      n3947, n5168, n3948, n5167, n3949, n5166, n5165, n5164, n5163, n5162, 
      n5161, n5160, n5089, n5088, n5087, n5086, n5085, n5084, n5083, n5082, 
      n5081, n5080, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, 
      n4008, n4009, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, 
      n4488, n4489, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, 
      n4568, n4569, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, 
      n4648, n4649, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, 
      n4728, n4729, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, 
      n4808, n4809, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n5199, 
      n3917, n5198, n3918, n5197, n3919, n5196, n5195, n5194, n5193, n5192, 
      n5191, n5190;

  EN210  g1( .A(n4777), .B(n4445), .Y(n4679) );
   AN210  g2( .A(A_2_port), .B(B_0_port), .Y(n4520) );
   BF003  g3( .A1(n4503), .A2(n3911), .B1(n5059), .B2(
                           n3912), .Y(n4678) );
   NA210  g4( .A(A_3_port), .B(B_0_port), .Y(n4273) );
   BF003  g5( .A1(n4502), .A2(n3909), .B1(n4114), .B2(
                           n3910), .Y(n4681) );
   NA210  g6( .A(A_4_port), .B(B_0_port), .Y(n4274) );
   BF003  g7( .A1(n4501), .A2(n4444), .B1(n4115), .B2(
                           n4447), .Y(n4227) );
   NA210  g8( .A(B_0_port), .B(A_5_port), .Y(n4275) );
   BF003  g9( .A1(n4500), .A2(n4442), .B1(n4116), .B2(
                           n4443), .Y(n5205) );
   NO210  g10( .A(n5103), .B(n4276), .Y(n4956) );
   EN210  g11( .A(n4960), .B(n4127), .Y(n4535) );
   EN2B0  g12( .A(n4185), .B(n4060), .Y(n4534) );
   EX2B0  g13( .A(n4186), .B(n4062), .Y(n4064) );
   EN2B0  g14( .A(n4188), .B(n4063), .Y(n4537) );
   BF003  g15( .A1(n4307), .A2(n4490), .B1(n4607), .B2(
                           n4065), .Y(n4489) );
   BF003  g16( .A1(n4306), .A2(n4491), .B1(n4608), .B2(
                           n4066), .Y(n4967) );
   EN210  g17( .A(n3942), .B(n4924), .Y(n4968) );
   EX2B0  g18( .A(n5145), .B(n4056), .Y(PRODUCT_6_port) );
   EX2B0  g19( .A(n4687), .B(n5066), .Y(PRODUCT_17_port) );
   EX210  g20( .A(n5147), .B(n5146), .Y(PRODUCT_14_port) );
   BF053  g21( .A1(n4546), .A2(n4226), .B1(n5165), .B2(
                           n5213), .Y(n5166) );
   IV110  g22( .A(B_13_port), .Y(n4811) );
   IV110  g23( .A(B_8_port), .Y(n4698) );
   IV110  g24( .A(A_13_port), .Y(n4285) );
   IV110  g25( .A(A_11_port), .Y(n4807) );
   IV110  g26( .A(B_5_port), .Y(n3873) );
   IV110  g27( .A(B_9_port), .Y(n4701) );
   NO210  g28( .A(n5064), .B(n4265), .Y(n4732) );
   NA410  g29( .A(n4640), .B(n5010), .C(n4733), .D(n4137), .Y(
                           n4731) );
   NA410  g30( .A(n4734), .B(n4731), .C(n4736), .D(n5082), .Y(
                           n4602) );
   BF053  g31( .A1(n3960), .A2(n3961), .B1(n5053), .B2(
                           n4329), .Y(n4865) );
   IV110  g32( .A(n4865), .Y(n4864) );
   BF053  g33( .A1(n5054), .A2(n4331), .B1(n5055), .B2(
                           n4862), .Y(n4863) );
   IV110  g34( .A(n4863), .Y(n4861) );
   BF053  g35( .A1(n4859), .A2(n3959), .B1(n5056), .B2(
                           n4335), .Y(n4860) );
   IV110  g36( .A(n4860), .Y(n4858) );
   BF053  g37( .A1(n4369), .A2(n3963), .B1(n5057), .B2(
                           n4338), .Y(n4857) );
   NO210  g38( .A(n5103), .B(n3873), .Y(n5036) );
   NO210  g39( .A(n3868), .B(n3871), .Y(n5035) );
   NA210  g40( .A(A_2_port), .B(B_3_port), .Y(n5038) );
   IV110  g41( .A(n4283), .Y(n4416) );
   IV110  g42( .A(n4712), .Y(n4417) );
   BF003  g43( .A1(n4936), .A2(n5072), .B1(n4275), .B2(
                           n4646), .Y(n4526) );
   BF003  g44( .A1(n4518), .A2(n5004), .B1(n4706), .B2(
                           n4568), .Y(n5005) );
   EN210  g45( .A(n4880), .B(n5005), .Y(n4883) );
   BF003  g46( .A1(n4517), .A2(n4565), .B1(n4702), .B2(
                           n4136), .Y(n4566) );
   BF003  g47( .A1(n4516), .A2(n4567), .B1(n5115), .B2(
                           n4564), .Y(n4882) );
   BF003  g48( .A1(n4515), .A2(n4134), .B1(n4699), .B2(
                           n4129), .Y(n4133) );
   IV110  g49( .A(n4726), .Y(n4585) );
   BF003  g50( .A1(n4514), .A2(n4135), .B1(n4703), .B2(
                           n4132), .Y(n4455) );
   EN210  g51( .A(n3971), .B(n3970), .Y(n3969) );
   EX210  g52( .A(n4379), .B(n3973), .Y(n3972) );
   EX2B0  g53( .A(n4521), .B(n4520), .Y(n4519) );
   EN210  g54( .A(n4382), .B(n4381), .Y(n4380) );
   EN210  g55( .A(n4096), .B(n4095), .Y(n4094) );
   EX2B0  g56( .A(n4913), .B(n4384), .Y(n4383) );
   EN210  g57( .A(n4093), .B(n4092), .Y(n4091) );
   EN210  g58( .A(n4387), .B(n4386), .Y(n4385) );
   EN210  g59( .A(n4090), .B(n4089), .Y(n4088) );
   EN210  g60( .A(n5031), .B(n4604), .Y(n4087) );
   BF003  g61( .A1(n3990), .A2(n4752), .B1(n4621), .B2(
                           n4753), .Y(n4336) );
   BF003  g62( .A1(n3989), .A2(n4332), .B1(n4622), .B2(
                           n4754), .Y(n4333) );
   BF053  g63( .A1(n4275), .A2(n5072), .B1(n4526), .B2(
                           n4094), .Y(n4153) );
   IV110  g64( .A(n4153), .Y(n4152) );
   BF053  g65( .A1(n5145), .A2(n4056), .B1(n4714), .B2(
                           n4152), .Y(n4151) );
   BF003  g66( .A1(n4715), .A2(n4151), .B1(n4804), .B2(
                           n4977), .Y(n4150) );
   BF053  g67( .A1(n4716), .A2(n4150), .B1(n5154), .B2(
                           n5153), .Y(n4149) );
   BF003  g68( .A1(n5105), .A2(n4980), .B1(n5125), .B2(
                           n4149), .Y(n4148) );
   BF003  g69( .A1(n5012), .A2(n4746), .B1(n4724), .B2(
                           n5166), .Y(n4433) );
   BF053  g70( .A1(n4055), .A2(n4054), .B1(n5126), .B2(
                           n4148), .Y(n4147) );
   BF053  g71( .A1(n4560), .A2(n4454), .B1(n4700), .B2(
                           n4131), .Y(n4559) );
   IV110  g72( .A(n4559), .Y(n4561) );
   BF053  g73( .A1(n4456), .A2(n4455), .B1(n4703), .B2(
                           n4135), .Y(n4562) );
   BF003  g74( .A1(n4416), .A2(n4761), .B1(n4283), .B2(
                           n4764), .Y(n5204) );
   IV110  g75( .A(n4562), .Y(n4563) );
   BF003  g76( .A1(n4415), .A2(n4229), .B1(n5132), .B2(
                           n4230), .Y(n4735) );
   BF053  g77( .A1(n4566), .A2(n4453), .B1(n4702), .B2(
                           n4565), .Y(n4564) );
   EX2B0  g78( .A(n4231), .B(n5133), .Y(n5160) );
   IV110  g79( .A(n4564), .Y(n4567) );
   BF003  g80( .A1(n4414), .A2(n4232), .B1(n5134), .B2(
                           n4233), .Y(n5182) );
   NA210  g81( .A(A_4_port), .B(B_12_port), .Y(n4191) );
   NA210  g82( .A(A_6_port), .B(B_10_port), .Y(n4192) );
   NA210  g83( .A(B_12_port), .B(A_11_port), .Y(n5139) );
   NA210  g84( .A(A_13_port), .B(B_10_port), .Y(n5140) );
   NA210  g85( .A(A_14_port), .B(B_9_port), .Y(n5141) );
   IV110  g86( .A(n4732), .Y(n4640) );
   IV110  g87( .A(n4279), .Y(n4835) );
   EX2B0  g88( .A(n4218), .B(n4871), .Y(n5148) );
   NO210  g89( .A(n5142), .B(n4484), .Y(n4384) );
   IV110  g90( .A(n4167), .Y(n4397) );
   IV110  g91( .A(n3883), .Y(n4836) );
   BF002  g92( .A1(n4600), .B1(n4053), .B2(n5007), .B3(
                           n4048), .Y(n4639) );
   NA210  g93( .A(B_9_port), .B(A_15_port), .Y(n5143) );
   IV110  g94( .A(n4203), .Y(n4817) );
   IV110  g95( .A(n3882), .Y(n3884) );
   NA210  g96( .A(n5065), .B(n4640), .Y(n4209) );
   IV110  g97( .A(n4202), .Y(n4818) );
   NA210  g98( .A(A_2_port), .B(B_14_port), .Y(n4041) );
   IV110  g99( .A(n4201), .Y(n4819) );
   NA210  g100( .A(n4367), .B(n4366), .Y(n4042) );
   BF053  g101( .A1(n5162), .A2(n4385), .B1(n4630), .B2(
                           n5163), .Y(n4631) );
   IV110  g102( .A(n4181), .Y(n4078) );
   IV110  g103( .A(n4180), .Y(n4079) );
   IV110  g104( .A(n4922), .Y(n4592) );
   IV110  g105( .A(n5123), .Y(n4081) );
   IV110  g106( .A(n3875), .Y(n3889) );
   IV110  g107( .A(n3874), .Y(n3890) );
   NO210  g108( .A(n4557), .B(n4392), .Y(n4944) );
   NA310  g109( .A(n4806), .B(n5007), .C(n4052), .Y(n4943) );
   BF056  g110( .A1(n5006), .A2(n4943), .B1(n4641), .B2(
                           n4944), .Y(n4394) );
   BF053  g111( .A1(n4191), .A2(n4237), .B1(n4469), .B2(
                           n4046), .Y(n4753) );
   IV110  g112( .A(n4753), .Y(n4752) );
   BF003  g113( .A1(n4618), .A2(n5184), .B1(n4750), .B2(
                           n3956), .Y(n4751) );
   BF003  g114( .A1(n4819), .A2(n4314), .B1(n4201), .B2(
                           n4315), .Y(n3967) );
   BF053  g115( .A1(n3957), .A2(n3958), .B1(n4619), .B2(
                           n5181), .Y(n4749) );
   EN210  g116( .A(n3966), .B(n4428), .Y(n3971) );
   IV110  g117( .A(n4749), .Y(n4748) );
   BF003  g118( .A1(n4818), .A2(n4316), .B1(n4202), .B2(
                           n4317), .Y(n3970) );
   BF053  g119( .A1(n3955), .A2(n3954), .B1(n4625), .B2(
                           n5177), .Y(n4747) );
   BF003  g120( .A1(n4817), .A2(n4318), .B1(n4203), .B2(
                           n4728), .Y(n3997) );
   NO210  g121( .A(n5104), .B(n4807), .Y(n5127) );
   IV110  g122( .A(B_7_port), .Y(n4276) );
   NA210  g123( .A(B_0_port), .B(A_10_port), .Y(n5126) );
   IV110  g124( .A(B_4_port), .Y(n3871) );
   NO210  g125( .A(n5104), .B(n5048), .Y(n5125) );
   IV110  g126( .A(B_15_port), .Y(n4142) );
   NA210  g127( .A(B_0_port), .B(A_8_port), .Y(n4716) );
   IV110  g128( .A(B_1_port), .Y(n5043) );
   NO210  g129( .A(n5104), .B(n4614), .Y(n4715) );
   IV110  g130( .A(B_6_port), .Y(n4277) );
   EX2B0  g131( .A(n4296), .B(n4016), .Y(n4013) );
   EN2B0  g132( .A(n4297), .B(n4014), .Y(n4011) );
   NA210  g133( .A(A_6_port), .B(B_8_port), .Y(n3882) );
   NA210  g134( .A(A_7_port), .B(B_7_port), .Y(n3883) );
   NA210  g135( .A(B_5_port), .B(A_9_port), .Y(n4279) );
   BF003  g136( .A1(n4399), .A2(n4838), .B1(n4549), .B2(
                           n4840), .Y(n4006) );
   NA210  g137( .A(B_4_port), .B(A_10_port), .Y(n4280) );
   EN210  g138( .A(n4550), .B(n4006), .Y(n4174) );
   NO210  g139( .A(n3870), .B(n4807), .Y(n4281) );
   BF003  g140( .A1(n3986), .A2(n4841), .B1(n4551), .B2(
                           n4842), .Y(n4173) );
   IV110  g141( .A(n4697), .Y(n4511) );
   IV110  g142( .A(n4129), .Y(n4134) );
   IV110  g143( .A(n4700), .Y(n4510) );
   IV110  g144( .A(n4703), .Y(n4514) );
   IV110  g145( .A(n4136), .Y(n4565) );
   EN210  g146( .A(n5206), .B(n5205), .Y(n4786) );
   BF053  g147( .A1(n4420), .A2(n4172), .B1(n4126), .B2(
                           n4421), .Y(n4049) );
   EN210  g148( .A(n4883), .B(n4882), .Y(n4881) );
   BF053  g149( .A1(n4549), .A2(n4838), .B1(n4550), .B2(
                           n4006), .Y(n4419) );
   EN210  g150( .A(n5209), .B(n5208), .Y(n5207) );
   IV110  g151( .A(n4419), .Y(n4005) );
   EN210  g152( .A(n4457), .B(n4877), .Y(n4880) );
   BF053  g153( .A1(n4551), .A2(n4841), .B1(n4174), .B2(
                           n4173), .Y(n4004) );
   EN210  g154( .A(n5212), .B(n5211), .Y(n5210) );
   IV110  g155( .A(n4004), .Y(n4003) );
   EN210  g156( .A(n4879), .B(n4878), .Y(n4877) );
   EN210  g157( .A(n4876), .B(n4458), .Y(n4457) );
   EN210  g158( .A(n4456), .B(n4455), .Y(n4454) );
   BF053  g159( .A1(n4615), .A2(n4155), .B1(n4031), .B2(
                           n4030), .Y(n5102) );
   EN210  g160( .A(n4025), .B(n4450), .Y(n4453) );
   IV110  g161( .A(n4658), .Y(n4237) );
   BF003  g162( .A1(n4576), .A2(n4952), .B1(n4207), .B2(
                           n4953), .Y(n4386) );
   BF053  g163( .A1(n4368), .A2(n4365), .B1(n4768), .B2(
                           n4767), .Y(n4236) );
   BF003  g164( .A1(n4826), .A2(n4950), .B1(n4208), .B2(
                           n4951), .Y(n4793) );
   BF053  g165( .A1(n4707), .A2(n3930), .B1(n4772), .B2(
                           n4771), .Y(n4235) );
   IV110  g166( .A(n4194), .Y(n4409) );
   EN210  g167( .A(n4680), .B(n4011), .Y(n4794) );
   IV110  g168( .A(n3894), .Y(n4846) );
   IV110  g169( .A(n4235), .Y(n4234) );
   IV110  g170( .A(n4193), .Y(n4410) );
   EX210  g171( .A(n4250), .B(n4010), .Y(n5215) );
   BF053  g172( .A1(n5070), .A2(n3897), .B1(n4117), .B2(
                           n4844), .Y(n4845) );
   BF053  g173( .A1(n4774), .A2(n4775), .B1(n4286), .B2(
                           n3925), .Y(n4233) );
   IV110  g174( .A(n4191), .Y(n4411) );
   EX2B0  g175( .A(n4949), .B(n4628), .Y(n4947) );
   IV110  g176( .A(n4845), .Y(n4843) );
   IV110  g177( .A(n4236), .Y(n4756) );
   IV110  g178( .A(n4189), .Y(n4413) );
   IV110  g179( .A(n5134), .Y(n4414) );
   IV110  g180( .A(n5132), .Y(n4415) );
   EN210  g181( .A(n4364), .B(n4363), .Y(n4362) );
   BF003  g182( .A1(n4184), .A2(n4059), .B1(n4061), .B2(
                           n4104), .Y(n4060) );
   EX210  g183( .A(n4361), .B(n4360), .Y(n4359) );
   BF053  g184( .A1(n4185), .A2(n4060), .B1(n4534), .B2(
                           n4535), .Y(n4062) );
   EN210  g185( .A(n3953), .B(n3952), .Y(n3951) );
   BF003  g186( .A1(n4581), .A2(n4850), .B1(n5139), .B2(
                           n4852), .Y(n4309) );
   BF003  g187( .A1(n4186), .A2(n4062), .B1(n4064), .B2(
                           n4105), .Y(n4063) );
   EN210  g188( .A(n4487), .B(n4309), .Y(n4909) );
   EN210  g189( .A(n3950), .B(n3949), .Y(n3948) );
   IV110  g190( .A(n4654), .Y(n4652) );
   BF053  g191( .A1(n4537), .A2(n4538), .B1(n4188), .B2(
                           n4063), .Y(n4065) );
   BF053  g192( .A1(n4112), .A2(n4650), .B1(n4111), .B2(
                           n4861), .Y(n4651) );
   EN210  g193( .A(n3947), .B(n3946), .Y(n3945) );
   IV110  g194( .A(n4651), .Y(n4649) );
   BF053  g195( .A1(n4607), .A2(n4490), .B1(n4489), .B2(
                           n4530), .Y(n4066) );
   BF053  g196( .A1(n4375), .A2(n4374), .B1(n4113), .B2(
                           n4864), .Y(n4648) );
   IV110  g197( .A(n4648), .Y(n4647) );
   BF053  g198( .A1(n4115), .A2(n4444), .B1(n4227), .B2(
                           n4786), .Y(n4228) );
   IV110  g199( .A(n4228), .Y(n4226) );
   BF053  g200( .A1(n4539), .A2(n4439), .B1(n4224), .B2(
                           n4783), .Y(n4225) );
   NA210  g201( .A(n4265), .B(n5064), .Y(n5065) );
   NO210  g202( .A(n5068), .B(n5067), .Y(n5066) );
   NA210  g203( .A(n4687), .B(n5066), .Y(n5009) );
   NO210  g204( .A(n5008), .B(n5009), .Y(n5010) );
   NA210  g205( .A(A_12_port), .B(B_13_port), .Y(n5069) );
   IV110  g206( .A(n4646), .Y(n5072) );
   BF053  g207( .A1(n5075), .A2(n4087), .B1(n4269), .B2(
                           n5074), .Y(n5073) );
   IV110  g208( .A(n5073), .Y(n5076) );
   IV110  g209( .A(n4119), .Y(n4405) );
   BF053  g210( .A1(n5031), .A2(n4604), .B1(n4606), .B2(
                           n4605), .Y(n5077) );
   EX210  g211( .A(n5148), .B(n4597), .Y(PRODUCT_30_port) );
   EX2B0  g212( .A(n5150), .B(n5149), .Y(PRODUCT_4_port) );
   EX210  g213( .A(n5152), .B(n5151), .Y(PRODUCT_12_port) );
   EX2B0  g214( .A(n4271), .B(n4272), .Y(PRODUCT_1_port) );
   EX2B0  g215( .A(n5154), .B(n5153), .Y(PRODUCT_8_port) );
   BF003  g216( .A1(n4210), .A2(n4209), .B1(n5010), .B2(
                           n4211), .Y(PRODUCT_19_port) );
   BF052  g217( .A1(n4213), .B1(n4212), .B2(n4168), .B3(
                           n4166), .Y(n4870) );
   EX210  g218( .A(n4031), .B(n4030), .Y(n4029) );
   EX2B0  g219( .A(n4028), .B(n4027), .Y(n4975) );
   EX210  g220( .A(n4974), .B(n4973), .Y(n4972) );
   NA210  g221( .A(n4632), .B(n5216), .Y(n4596) );
   NA311  g222( .A(n4398), .B(n4988), .C(n4596), .Y(n4730) );
   BF056  g223( .A1(n4730), .A2(n4990), .B1(n4168), .B2(
                           n4212), .Y(n4694) );
   BF053  g224( .A1(n4726), .A2(n4432), .B1(n4729), .B2(
                           n4910), .Y(n4558) );
   BF053  g225( .A1(n4727), .A2(n4907), .B1(n5140), .B2(
                           n4853), .Y(n4728) );
   IV110  g226( .A(n4728), .Y(n4318) );
   BF053  g227( .A1(n4908), .A2(n4909), .B1(n5135), .B2(
                           n4435), .Y(n4317) );
   NA210  g228( .A(A_8_port), .B(B_12_port), .Y(n4543) );
   NA210  g229( .A(B_11_port), .B(A_9_port), .Y(n4544) );
   NA210  g230( .A(A_14_port), .B(B_7_port), .Y(n4545) );
   NA210  g231( .A(n5033), .B(n5032), .Y(n5039) );
   NA210  g232( .A(B_2_port), .B(A_0_port), .Y(n4523) );
   NA210  g233( .A(A_1_port), .B(B_1_port), .Y(n4524) );
   NA210  g234( .A(A_2_port), .B(B_1_port), .Y(n4089) );
   OR210  g235( .A(n4523), .B(n4524), .Y(n4090) );
   NA210  g236( .A(A_3_port), .B(B_1_port), .Y(n4269) );
   NA210  g237( .A(A_4_port), .B(B_1_port), .Y(n4270) );
   NO210  g238( .A(n5043), .B(n4187), .Y(n5042) );
   NA210  g239( .A(B_1_port), .B(A_6_port), .Y(n5044) );
   NO210  g240( .A(n5043), .B(n4614), .Y(n5045) );
   IV110  g241( .A(n4205), .Y(n4578) );
   EN210  g242( .A(n4453), .B(n4566), .Y(n4456) );
   IV110  g243( .A(n4206), .Y(n4577) );
   BF003  g244( .A1(n4513), .A2(n4563), .B1(n5116), .B2(
                           n4562), .Y(n4999) );
   IV110  g245( .A(n4207), .Y(n4576) );
   EN210  g246( .A(n4881), .B(n4999), .Y(n4532) );
   IV110  g247( .A(n4208), .Y(n4826) );
   IV110  g248( .A(n4212), .Y(n4988) );
   IV110  g249( .A(n4946), .Y(n5163) );
   IV110  g250( .A(n5159), .Y(n5158) );
   EN210  g251( .A(n5034), .B(n5037), .Y(n5040) );
   EN210  g252( .A(n5039), .B(n5038), .Y(n5037) );
   EN210  g253( .A(n5036), .B(n5035), .Y(n5034) );
   EN210  g254( .A(n5033), .B(n5032), .Y(n5031) );
   NO210  g255( .A(n5103), .B(n4277), .Y(n4017) );
   EN210  g256( .A(n4606), .B(n4605), .Y(n4604) );
   NA210  g257( .A(A_2_port), .B(B_5_port), .Y(n4958) );
   NA210  g258( .A(n4965), .B(n4017), .Y(n4959) );
   EN210  g259( .A(n4780), .B(n4219), .Y(n4785) );
   NA210  g260( .A(A_2_port), .B(B_4_port), .Y(n4962) );
   IV110  g261( .A(n4110), .Y(n4506) );
   IV110  g262( .A(n4109), .Y(n4507) );
   IV110  g263( .A(n4115), .Y(n4501) );
   IV110  g264( .A(n4116), .Y(n4500) );
   IV110  g265( .A(n4539), .Y(n4499) );
   BF003  g266( .A1(n4305), .A2(n4493), .B1(n4609), .B2(
                           n4492), .Y(n5029) );
   EN210  g267( .A(n4101), .B(n5029), .Y(n4971) );
   EN210  g268( .A(n4105), .B(n4064), .Y(n4028) );
   EN210  g269( .A(n4104), .B(n4061), .Y(n4974) );
   BF003  g270( .A1(n4304), .A2(n4160), .B1(n4610), .B2(
                           n4163), .Y(n4973) );
   BF053  g271( .A1(n4452), .A2(n4451), .B1(n4450), .B2(
                           n4025), .Y(n4568) );
   BF003  g272( .A1(n4413), .A2(n4234), .B1(n4189), .B2(
                           n4235), .Y(n5178) );
   BF003  g273( .A1(n4412), .A2(n4756), .B1(n4190), .B2(
                           n4236), .Y(n5175) );
   EN210  g274( .A(n4043), .B(n5175), .Y(n4469) );
   BF003  g275( .A1(n4411), .A2(n4237), .B1(n4191), .B2(
                           n4658), .Y(n4046) );
   EN210  g276( .A(n4045), .B(n5178), .Y(n4472) );
   EN2B0  g277( .A(n4192), .B(n4660), .Y(n4471) );
   IV110  g278( .A(n4242), .Y(n4240) );
   BF053  g279( .A1(n4270), .A2(n5076), .B1(n4096), .B2(
                           n4095), .Y(n4239) );
   BF003  g280( .A1(n5042), .A2(n4239), .B1(n5193), .B2(
                           n4972), .Y(n5194) );
   NA210  g281( .A(A_12_port), .B(B_12_port), .Y(n5144) );
   IV110  g282( .A(n3881), .Y(n3885) );
   NA210  g283( .A(A_10_port), .B(B_14_port), .Y(n4199) );
   IV110  g284( .A(n4245), .Y(n3931) );
   NA210  g285( .A(A_9_port), .B(B_15_port), .Y(n4200) );
   IV110  g286( .A(n4199), .Y(n4820) );
   IV110  g287( .A(n3878), .Y(n3887) );
   NA210  g288( .A(n4267), .B(n4635), .Y(n5082) );
   NA210  g289( .A(A_11_port), .B(B_13_port), .Y(n4201) );
   IV110  g290( .A(n5144), .Y(n4821) );
   IV110  g291( .A(n3877), .Y(n3888) );
   NA210  g292( .A(n4800), .B(n4050), .Y(n4570) );
   NA210  g293( .A(A_13_port), .B(B_11_port), .Y(n4202) );
   IV110  g294( .A(n5143), .Y(n4822) );
   IV110  g295( .A(n4765), .Y(n4762) );
   IV110  g296( .A(n4869), .Y(n4166) );
   IV110  g297( .A(n5070), .Y(n4407) );
   EN210  g298( .A(n4359), .B(n4759), .Y(n4364) );
   EN210  g299( .A(n4282), .B(n5096), .Y(n4363) );
   BF003  g300( .A1(n4833), .A2(n4762), .B1(n3876), .B2(
                           n4765), .Y(n4763) );
   NA410  g301( .A(n4596), .B(n4869), .C(n4602), .D(n4988), .Y(
                           n4213) );
   BF053  g302( .A1(n3974), .A2(n3975), .B1(n4553), .B2(
                           n4003), .Y(n4798) );
   BF053  g303( .A1(n4555), .A2(n4942), .B1(n4554), .B2(
                           n4005), .Y(n4875) );
   IV110  g304( .A(n4293), .Y(n5019) );
   NO210  g305( .A(n4050), .B(n4800), .Y(n4216) );
   IV110  g306( .A(n4724), .Y(n5012) );
   OR310  g307( .A(n4986), .B(n4051), .C(n4398), .Y(n4215) );
   IV110  g308( .A(n4723), .Y(n5013) );
   NA410  g309( .A(n4571), .B(n4048), .C(n5007), .D(n4053), .Y(
                           n4217) );
   IV110  g310( .A(n4722), .Y(n5014) );
   IV110  g311( .A(n4747), .Y(n4338) );
   EN210  g312( .A(n3969), .B(n3997), .Y(n4379) );
   EX2B0  g313( .A(n3972), .B(n4558), .Y(n4381) );
   BF003  g314( .A1(n4408), .A2(n3895), .B1(n5069), .B2(
                           n3896), .Y(n5107) );
   BF003  g315( .A1(n4407), .A2(n3897), .B1(n5070), .B2(
                           n3899), .Y(n4844) );
   EN210  g316( .A(n4117), .B(n4844), .Y(n5108) );
   BF003  g317( .A1(n4406), .A2(n4427), .B1(n4118), .B2(
                           n4837), .Y(n4425) );
   IV110  g318( .A(n3910), .Y(n3909) );
   BF053  g319( .A1(n4114), .A2(n3909), .B1(n4682), .B2(
                           n4681), .Y(n3908) );
   IV110  g320( .A(n3908), .Y(n3907) );
   EX210  g321( .A(n4964), .B(n4961), .Y(n4104) );
   IV110  g322( .A(n5025), .Y(n5024) );
   BF053  g323( .A1(n5022), .A2(n4357), .B1(n4181), .B2(
                           n4917), .Y(n5023) );
   EN210  g324( .A(n4623), .B(n4333), .Y(n4904) );
   IV110  g325( .A(n5023), .Y(n5021) );
   BF003  g326( .A1(n3988), .A2(n4755), .B1(n4624), .B2(
                           n5176), .Y(n4903) );
   BF053  g327( .A1(n4097), .A2(n4358), .B1(n4180), .B2(
                           n4921), .Y(n4595) );
   EN210  g328( .A(n4902), .B(n4336), .Y(n3955) );
   IV110  g329( .A(n4595), .Y(n4594) );
   BF003  g330( .A1(n3987), .A2(n5177), .B1(n4625), .B2(
                           n5179), .Y(n3954) );
   BF003  g331( .A1(n3886), .A2(n3931), .B1(n3880), .B2(n4245),
                           .Y(n3932) );
   BF003  g332( .A1(n3887), .A2(n4243), .B1(n3878), .B2(n4244),
                           .Y(n3926) );
   BF003  g333( .A1(n3888), .A2(n4240), .B1(n3877), .B2(n4242),
                           .Y(n3952) );
   EN2B0  g334( .A(n4808), .B(n5185), .Y(n4038) );
   EN210  g335( .A(n4887), .B(n5095), .Y(n4039) );
   BF003  g336( .A1(n3889), .A2(n5028), .B1(n3875), .B2(n5030),
                           .Y(n4888) );
   EN210  g337( .A(n4467), .B(n4676), .Y(n4889) );
   NA210  g338( .A(B_0_port), .B(A_6_port), .Y(n4714) );
   NA210  g339( .A(B_3_port), .B(A_12_port), .Y(n4713) );
   NA210  g340( .A(B_4_port), .B(A_11_port), .Y(n4712) );
   NO210  g341( .A(n5103), .B(n5124), .Y(n4355) );
   NA210  g342( .A(n3937), .B(n3936), .Y(n4352) );
   NA210  g343( .A(A_2_port), .B(B_10_port), .Y(n4351) );
   NA210  g344( .A(B_4_port), .B(A_8_port), .Y(n5123) );
   NA210  g345( .A(B_5_port), .B(A_6_port), .Y(n5122) );
   NA210  g350( .A(A_5_port), .B(B_6_port), .Y(n5121) );
   NA210  g351( .A(A_4_port), .B(B_7_port), .Y(n5120) );
   NA210  g352( .A(B_2_port), .B(A_12_port), .Y(n4282) );
   EX210  g353( .A(n4172), .B(n4420), .Y(n4177) );
   NA210  g354( .A(B_1_port), .B(A_14_port), .Y(n4283) );
   EN210  g355( .A(n4169), .B(n4552), .Y(n4391) );
   NO210  g356( .A(n3869), .B(n4285), .Y(n4284) );
   EX2B0  g357( .A(n5109), .B(n4945), .Y(n3980) );
   NA210  g358( .A(A_6_port), .B(B_9_port), .Y(n4286) );
   BF003  g359( .A1(n3985), .A2(n4003), .B1(n4553), .B2(
                           n4004), .Y(n3974) );
   NO210  g360( .A(n4187), .B(n4705), .Y(n4287) );
   BF003  g361( .A1(n4005), .A2(n3984), .B1(n4419), .B2(
                           n4554), .Y(n4942) );
   BF053  g362( .A1(n3971), .A2(n3970), .B1(n4202), .B2(
                           n4316), .Y(n4002) );
   IV110  g363( .A(n3919), .Y(n4446) );
   IV110  g364( .A(n4002), .Y(n4001) );
   IV110  g365( .A(n4107), .Y(n4926) );
   BF053  g366( .A1(n4119), .A2(n4001), .B1(n5111), .B2(
                           n5110), .Y(n4000) );
   BF053  g367( .A1(n5099), .A2(n4966), .B1(n4616), .B2(
                           n5100), .Y(n5101) );
   IV110  g368( .A(n4108), .Y(n4508) );
   EN210  g369( .A(n4452), .B(n4451), .Y(n4450) );
   IV110  g370( .A(n4000), .Y(n3999) );
   IV110  g371( .A(n5101), .Y(n5098) );
   IV110  g372( .A(n4113), .Y(n4504) );
   EN210  g373( .A(n4449), .B(n4026), .Y(n4025) );
   BF053  g374( .A1(n4170), .A2(n4171), .B1(n4121), .B2(
                           n3999), .Y(n4176) );
   BF053  g375( .A1(n5041), .A2(n5098), .B1(n4971), .B2(
                           n4970), .Y(n5097) );
   IV110  g376( .A(n4111), .Y(n4505) );
   EN210  g377( .A(n4018), .B(n4021), .Y(n4024) );
   BF003  g378( .A1(n4809), .A2(n5097), .B1(n5095), .B2(
                           n4887), .Y(n5096) );
   BF053  g379( .A1(n3875), .A2(n5028), .B1(n4889), .B2(
                           n4888), .Y(n5094) );
   BF003  g380( .A1(n4927), .A2(n4446), .B1(n5060), .B2(
                           n3919), .Y(n4445) );
   BF053  g381( .A1(n4676), .A2(n4467), .B1(n3874), .B2(
                           n5026), .Y(n5093) );
   EN2B0  g382( .A(n4629), .B(n4948), .Y(n5164) );
   BF003  g383( .A1(n4825), .A2(n5163), .B1(n4630), .B2(
                           n4946), .Y(n5162) );
   EN210  g384( .A(n4792), .B(n4631), .Y(n4263) );
   EN210  g385( .A(n4388), .B(n4947), .Y(n3860) );
   EN2B0  g386( .A(n4633), .B(n5161), .Y(n3859) );
   IV110  g387( .A(n4619), .Y(n3992) );
   IV110  g388( .A(n5166), .Y(n4746) );
   IV110  g389( .A(n5180), .Y(n3922) );
   BF053  g390( .A1(n4293), .A2(n5167), .B1(n4249), .B2(
                           n5214), .Y(n4745) );
   BF003  g391( .A1(n4083), .A2(n5000), .B1(n5122), .B2(
                           n4998), .Y(n3943) );
   IV110  g392( .A(n4745), .Y(n4744) );
   BF003  g393( .A1(n4082), .A2(n4997), .B1(n5117), .B2(
                           n4996), .Y(n4924) );
   BF053  g394( .A1(n4292), .A2(n4221), .B1(n5212), .B2(
                           n5211), .Y(n4743) );
   BF003  g395( .A1(n4081), .A2(n4925), .B1(n5123), .B2(
                           n4923), .Y(n4102) );
   IV110  g396( .A(n4743), .Y(n4742) );
   BF003  g397( .A1(n4080), .A2(n4592), .B1(n4179), .B2(
                           n4922), .Y(n4591) );
   EN210  g398( .A(n4356), .B(n4591), .Y(n4097) );
   BF003  g399( .A1(n4079), .A2(n4921), .B1(n4180), .B2(
                           n4918), .Y(n4358) );
   BF003  g400( .A1(n4078), .A2(n4917), .B1(n4181), .B2(
                           n4916), .Y(n5022) );
   EN210  g401( .A(n4357), .B(n5022), .Y(n4100) );
   IV110  g402( .A(n4066), .Y(n4491) );
   EN210  g403( .A(n4899), .B(n4735), .Y(n5067) );
   BF053  g404( .A1(n4968), .A2(n4967), .B1(n4608), .B2(
                           n4491), .Y(n4492) );
   EN2B0  g405( .A(n4362), .B(n4763), .Y(n5146) );
   IV110  g406( .A(n4492), .Y(n4493) );
   IV110  g407( .A(n4225), .Y(n4223) );
   EN210  g408( .A(n4969), .B(n4766), .Y(n5151) );
   BF053  g409( .A1(n4785), .A2(n4784), .B1(n4544), .B2(
                           n4655), .Y(n4222) );
   BF053  g410( .A1(n4349), .A2(n3943), .B1(n5122), .B2(
                           n5000), .Y(n4494) );
   BF003  g411( .A1(n5160), .A2(n4896), .B1(n5133), .B2(
                           n4231), .Y(n5161) );
   EN2B0  g412( .A(n4029), .B(n5187), .Y(n4054) );
   BF053  g413( .A1(n4633), .A2(n5161), .B1(n3859), .B2(
                           n3860), .Y(n5159) );
   IV110  g414( .A(n4494), .Y(n4495) );
   BF053  g415( .A1(n3863), .A2(n3862), .B1(n4634), .B2(
                           n5158), .Y(n4261) );
   EN210  g416( .A(n4972), .B(n5193), .Y(n4056) );
   BF053  g417( .A1(n4198), .A2(n5091), .B1(n4901), .B2(
                           n4900), .Y(n5157) );
   BF053  g418( .A1(n5155), .A2(n3858), .B1(n4636), .B2(
                           n5156), .Y(n5061) );
   NO210  g419( .A(n4574), .B(n4573), .Y(n4572) );
   OR210  g420( .A(n4635), .B(n4267), .Y(n4137) );
   NA210  g421( .A(n4571), .B(n4570), .Y(n4569) );
   IV110  g422( .A(n4121), .Y(n4404) );
   BF053  g423( .A1(n4964), .A2(n4961), .B1(n4963), .B2(
                           n4962), .Y(n5078) );
   IV110  g424( .A(n4053), .Y(n4574) );
   BF053  g425( .A1(n4127), .A2(n4960), .B1(n4278), .B2(
                           n5080), .Y(n5079) );
   IV110  g426( .A(n4944), .Y(n5007) );
   NO210  g427( .A(n3869), .B(n3868), .Y(n4092) );
   IV110  g428( .A(n5079), .Y(n4128) );
   NO210  g429( .A(n3870), .B(n5103), .Y(n4093) );
   IV110  g430( .A(n4216), .Y(n4571) );
   NA210  g431( .A(B_2_port), .B(A_2_port), .Y(n4605) );
   BF053  g432( .A1(n4957), .A2(n4527), .B1(n4959), .B2(
                           n4958), .Y(n4129) );
   NA210  g433( .A(n4092), .B(n4093), .Y(n4606) );
   IV110  g434( .A(n3965), .Y(n4915) );
   NO210  g435( .A(n3870), .B(n3868), .Y(n5033) );
   BF053  g436( .A1(n4106), .A2(n4529), .B1(n4697), .B2(
                           n4128), .Y(n4130) );
   NO210  g437( .A(n5103), .B(n3871), .Y(n5032) );
   NA210  g438( .A(B_2_port), .B(A_3_port), .Y(n3872) );
   NA210  g439( .A(B_3_port), .B(A_7_port), .Y(n4607) );
   NA210  g440( .A(B_3_port), .B(A_8_port), .Y(n4608) );
   NA210  g441( .A(B_3_port), .B(A_9_port), .Y(n4609) );
   EX210  g442( .A(n4971), .B(n4970), .Y(n4969) );
   EN210  g443( .A(n4968), .B(n4967), .Y(n4966) );
   EX210  g444( .A(n4538), .B(n4537), .Y(n4536) );
   IV110  g445( .A(n5030), .Y(n5028) );
   EX210  g446( .A(n4535), .B(n4534), .Y(n4533) );
   BF053  g447( .A1(n4102), .A2(n4103), .B1(n5123), .B2(
                           n4925), .Y(n5027) );
   EN210  g448( .A(n4532), .B(n4531), .Y(n4530) );
   IV110  g449( .A(n5027), .Y(n5026) );
   EX210  g450( .A(n4529), .B(n4106), .Y(n4105) );
   BF053  g451( .A1(n4100), .A2(n4099), .B1(n4182), .B2(
                           n4498), .Y(n5025) );
   NA210  g452( .A(A_13_port), .B(B_8_port), .Y(n4546) );
   NA210  g453( .A(B_10_port), .B(A_11_port), .Y(n4547) );
   NA210  g454( .A(A_7_port), .B(B_14_port), .Y(n4548) );
   NA210  g455( .A(A_6_port), .B(B_15_port), .Y(n4289) );
   NA210  g456( .A(A_8_port), .B(B_13_port), .Y(n4290) );
   NA210  g457( .A(B_12_port), .B(A_9_port), .Y(n4291) );
   NA210  g458( .A(B_11_port), .B(A_10_port), .Y(n4292) );
   NA210  g459( .A(B_12_port), .B(A_15_port), .Y(n4126) );
   BF003  g460( .A1(n3890), .A2(n5026), .B1(n3874), .B2(n5027
                           ), .Y(n4676) );
   NA210  g461( .A(A_13_port), .B(B_14_port), .Y(n4549) );
   EN210  g462( .A(n4464), .B(n4241), .Y(n4886) );
   NA210  g463( .A(A_12_port), .B(B_15_port), .Y(n4550) );
   BF003  g464( .A1(n3891), .A2(n5024), .B1(n4816), .B2(n5025
                           ), .Y(n4241) );
   IV110  g465( .A(n5135), .Y(n4584) );
   IV110  g466( .A(n5136), .Y(n4583) );
   IV110  g467( .A(n5137), .Y(n4582) );
   IV110  g468( .A(n5139), .Y(n4581) );
   IV110  g469( .A(n5140), .Y(n4580) );
   NA210  g470( .A(B_1_port), .B(A_8_port), .Y(n5046) );
   IV110  g471( .A(n5141), .Y(n4579) );
   NO210  g472( .A(n5043), .B(n5048), .Y(n5047) );
   BF003  g473( .A1(n4937), .A2(n5071), .B1(n4274), .B2(n4644
                           ), .Y(n5150) );
   NA210  g474( .A(B_1_port), .B(A_10_port), .Y(n5049) );
   NO210  g475( .A(n5043), .B(n4807), .Y(n5050) );
   NA210  g476( .A(B_1_port), .B(A_12_port), .Y(n4808) );
   NO210  g477( .A(n3869), .B(n4807), .Y(n4809) );
   NA210  g478( .A(B_5_port), .B(A_8_port), .Y(n4810) );
   NA210  g479( .A(A_5_port), .B(B_12_port), .Y(n4621) );
   NA210  g480( .A(A_3_port), .B(B_14_port), .Y(n4622) );
   NA210  g481( .A(A_2_port), .B(B_15_port), .Y(n4623) );
   IV110  g482( .A(n5157), .Y(n5156) );
   IV110  g483( .A(n4140), .Y(n4733) );
   EN210  g484( .A(n3944), .B(n3932), .Y(n3947) );
   BF003  g485( .A1(n3885), .A2(n4246), .B1(n3881), .B2(
                           n4667), .Y(n3946) );
   EN210  g486( .A(n3945), .B(n3926), .Y(n3950) );
   BF003  g487( .A1(n3884), .A2(n4668), .B1(n3882), .B2(
                           n4670), .Y(n3949) );
   BF003  g488( .A1(n4836), .A2(n4671), .B1(n3883), .B2(
                           n4672), .Y(n4342) );
   EN210  g489( .A(n3948), .B(n4342), .Y(n3953) );
   BF003  g490( .A1(n4835), .A2(n4673), .B1(n4279), .B2(
                           n4674), .Y(n4347) );
   EN210  g491( .A(n3951), .B(n4347), .Y(n4361) );
   BF003  g492( .A1(n4073), .A2(n4655), .B1(n4544), .B2(
                           n4656), .Y(n4784) );
   NA210  g493( .A(n5036), .B(n5035), .Y(n4963) );
   EN210  g494( .A(n4783), .B(n4224), .Y(n5206) );
   NA210  g495( .A(A_3_port), .B(B_4_port), .Y(n4278) );
   EN210  g496( .A(n4786), .B(n4227), .Y(n4682) );
   IV110  g497( .A(n5116), .Y(n4513) );
   NA210  g498( .A(B_4_port), .B(A_4_port), .Y(n4697) );
   IV110  g499( .A(n4009), .Y(n4007) );
   BF003  g500( .A1(n4072), .A2(n3907), .B1(n4545), .B2(
                           n3908), .Y(n4251) );
   IV110  g501( .A(n5115), .Y(n4516) );
   NO210  g502( .A(n5103), .B(n4698), .Y(n4020) );
   BF053  g503( .A1(n4205), .A2(n4007), .B1(n4787), .B2(
                           n4788), .Y(n4955) );
   BF003  g504( .A1(n4071), .A2(n4226), .B1(n4546), .B2(
                           n4228), .Y(n5165) );
   IV110  g505( .A(n4568), .Y(n5004) );
   NO210  g506( .A(n3868), .B(n4276), .Y(n4019) );
   IV110  g507( .A(n4955), .Y(n4954) );
   IV110  g508( .A(n5117), .Y(n4082) );
   IV110  g509( .A(n5122), .Y(n4083) );
   IV110  g510( .A(n5121), .Y(n4084) );
   IV110  g511( .A(n5120), .Y(n4085) );
   EX210  g512( .A(n4611), .B(n4159), .Y(n4157) );
   EN210  g513( .A(n4612), .B(n4158), .Y(n4027) );
   EX210  g514( .A(n4613), .B(n4156), .Y(n4154) );
   EN210  g515( .A(n4615), .B(n4155), .Y(n4030) );
   EN210  g516( .A(n4530), .B(n4489), .Y(n4031) );
   EN210  g517( .A(n4469), .B(n4046), .Y(n4045) );
   EN210  g518( .A(n4472), .B(n4471), .Y(n4470) );
   EN210  g519( .A(n4475), .B(n4474), .Y(n4473) );
   EN210  g520( .A(n4478), .B(n4477), .Y(n4476) );
   EX210  g521( .A(n4898), .B(n4897), .Y(n4896) );
   BF053  g522( .A1(n4978), .A2(n4979), .B1(n5044), .B2(
                           n5194), .Y(n5192) );
   BF003  g523( .A1(n5190), .A2(n4975), .B1(n5045), .B2(
                           n5192), .Y(n5191) );
   BF053  g524( .A1(n5046), .A2(n5191), .B1(n4981), .B2(
                           n4982), .Y(n5189) );
   BF003  g525( .A1(n5047), .A2(n5189), .B1(n5187), .B2(
                           n4029), .Y(n5188) );
   BF053  g526( .A1(n5049), .A2(n5188), .B1(n4984), .B2(
                           n4985), .Y(n5186) );
   BF003  g527( .A1(n5050), .A2(n5186), .B1(n4766), .B2(
                           n4969), .Y(n5185) );
   BF053  g528( .A1(n4808), .A2(n5185), .B1(n4038), .B2(
                           n4039), .Y(n4765) );
   EX2B0  g529( .A(n4601), .B(n3865), .Y(PRODUCT_23_port) );
   EX2B0  g530( .A(n4138), .B(n3866), .Y(PRODUCT_20_port) );
   EX2B0  g531( .A(n4575), .B(n3867), .Y(PRODUCT_27_port) );
   EX210  g532( .A(n3924), .B(n4284), .Y(n5090) );
   BF003  g533( .A1(n4832), .A2(n3925), .B1(n4286), .B2(
                           n3927), .Y(n4774) );
   EX2B0  g534( .A(n3928), .B(n4287), .Y(n4659) );
   BF003  g535( .A1(n4831), .A2(n4238), .B1(n4288), .B2(
                           n3929), .Y(n4657) );
   EN210  g536( .A(n4769), .B(n4657), .Y(n4772) );
   BF003  g537( .A1(n4830), .A2(n3930), .B1(n4707), .B2(
                           n3933), .Y(n4771) );
   EN210  g538( .A(n4770), .B(n4659), .Y(n4775) );
   EX210  g539( .A(n4268), .B(n4795), .Y(n4267) );
   BF003  g540( .A1(n4689), .A2(n4688), .B1(n4691), .B2(
                           n4690), .Y(n4687) );
   EN2B0  g541( .A(n4693), .B(n4692), .Y(n5008) );
   NA410  g542( .A(n4052), .B(n5007), .C(n4806), .D(n4053), .Y(
                           n4941) );
   IV110  g543( .A(n4721), .Y(n5015) );
   IV110  g544( .A(n4719), .Y(n5016) );
   IV110  g545( .A(n4718), .Y(n5017) );
   IV110  g546( .A(n4717), .Y(n5018) );
   IV110  g547( .A(n4617), .Y(n4929) );
   IV110  g548( .A(n4626), .Y(n4928) );
   EN2B0  g549( .A(n5049), .B(n5188), .Y(n4984) );
   EX210  g550( .A(n5050), .B(n5186), .Y(n4766) );
   EX210  g551( .A(n5097), .B(n4809), .Y(n5095) );
   BF053  g552( .A1(n4251), .A2(n4252), .B1(n4545), .B2(
                           n3907), .Y(n3906) );
   IV110  g553( .A(n3906), .Y(n3905) );
   BF053  g554( .A1(n4486), .A2(n4485), .B1(n4725), .B2(
                           n3905), .Y(n4914) );
   IV110  g555( .A(n4630), .Y(n4825) );
   BF053  g556( .A1(n4723), .A2(n4744), .B1(n4483), .B2(
                           n4482), .Y(n3904) );
   IV110  g557( .A(n4603), .Y(n4168) );
   IV110  g558( .A(n3904), .Y(n4856) );
   IV110  g559( .A(n4634), .Y(n4824) );
   BF053  g560( .A1(n4854), .A2(n4686), .B1(n4717), .B2(
                           n4323), .Y(n4855) );
   IV110  g561( .A(n4636), .Y(n4823) );
   BF053  g562( .A1(n4591), .A2(n4356), .B1(n4179), .B2(
                           n4592), .Y(n4593) );
   EN210  g563( .A(n4905), .B(n3921), .Y(n3958) );
   EX2B0  g564( .A(n4618), .B(n5184), .Y(n4750) );
   EN2B0  g565( .A(n5051), .B(n4751), .Y(n3918) );
   BF003  g566( .A1(n4935), .A2(n4748), .B1(n5052), .B2(
                           n4749), .Y(n4371) );
   BF003  g567( .A1(n4934), .A2(n4329), .B1(n5053), .B2(
                           n4330), .Y(n3960) );
   BF003  g568( .A1(n4331), .A2(n4933), .B1(n4334), .B2(
                           n5054), .Y(n4862) );
   BF053  g569( .A1(n5147), .A2(n5146), .B1(n5130), .B2(
                           n4144), .Y(n5092) );
   BF003  g570( .A1(n5131), .A2(n5092), .B1(n3864), .B2(
                           n5203), .Y(n5068) );
   BF003  g571( .A1(n5090), .A2(n5200), .B1(n4284), .B2(
                           n3924), .Y(n5091) );
   NA210  g572( .A(A_3_port), .B(B_8_port), .Y(n5119) );
   NO210  g573( .A(n3868), .B(n4705), .Y(n3936) );
   NO210  g574( .A(n5103), .B(n5118), .Y(n3937) );
   EX2B0  g575( .A(n4572), .B(n4394), .Y(PRODUCT_28_port) );
   EX2B0  g576( .A(n4393), .B(n4175), .Y(n4392) );
   EN210  g577( .A(n4391), .B(n4390), .Y(n4389) );
   EN210  g578( .A(n3983), .B(n3979), .Y(n3982) );
   EN210  g579( .A(n3981), .B(n3980), .Y(n3979) );
   EN210  g580( .A(n3978), .B(n3977), .Y(n3976) );
   EX210  g581( .A(n3975), .B(n3974), .Y(n4178) );
   EN210  g582( .A(n4555), .B(n4942), .Y(n3975) );
   EN210  g583( .A(n4178), .B(n4049), .Y(n3978) );
   BF053  g584( .A1(n4478), .A2(n4477), .B1(n4195), .B2(
                           n4666), .Y(n4431) );
   BF003  g585( .A1(n4294), .A2(n4431), .B1(n4429), .B2(
                           n4253), .Y(n4430) );
   BF053  g586( .A1(n4295), .A2(n4430), .B1(n4015), .B2(
                           n4256), .Y(n4016) );
   BF003  g587( .A1(n4013), .A2(n4677), .B1(n4296), .B2(
                           n4016), .Y(n4014) );
   BF053  g588( .A1(n4011), .A2(n4680), .B1(n4297), .B2(
                           n4014), .Y(n4012) );
   BF003  g589( .A1(n4298), .A2(n4012), .B1(n4010), .B2(
                           n4250), .Y(n5142) );
   IV110  g590( .A(n4704), .Y(n4509) );
   BF053  g591( .A1(n4008), .A2(n4476), .B1(n4196), .B2(
                           n5085), .Y(n4009) );
   BF003  g592( .A1(n4926), .A2(n3916), .B1(n4107), .B2(
                           n3917), .Y(n4778) );
   IV110  g593( .A(n5093), .Y(n4675) );
   BF003  g594( .A1(n4508), .A2(n4866), .B1(n4108), .B2(
                           n3915), .Y(n4440) );
   BF053  g595( .A1(n4468), .A2(n4886), .B1(n4810), .B2(
                           n4586), .Y(n4674) );
   BF003  g596( .A1(n4507), .A2(n4448), .B1(n4109), .B2(
                           n4857), .Y(n4377) );
   IV110  g597( .A(n4674), .Y(n4673) );
   BF003  g598( .A1(n4506), .A2(n4858), .B1(n4110), .B2(
                           n4860), .Y(n4653) );
   BF003  g599( .A1(n4505), .A2(n4861), .B1(n4111), .B2(
                           n4863), .Y(n4650) );
   EN210  g600( .A(n4112), .B(n4650), .Y(n4375) );
   BF003  g601( .A1(n4504), .A2(n4864), .B1(n4113), .B2(
                           n4865), .Y(n4374) );
   BF053  g602( .A1(n5209), .A2(n5208), .B1(n4290), .B2(
                           n5172), .Y(n4741) );
   IV110  g603( .A(B_10_port), .Y(n4705) );
   IV110  g604( .A(n4741), .Y(n4740) );
   IV110  g605( .A(n3872), .Y(n4940) );
   BF053  g606( .A1(n4548), .A2(n5169), .B1(n4289), .B2(
                           n4738), .Y(n4739) );
   BF003  g607( .A1(n4077), .A2(n4498), .B1(n4182), .B2(
                           n4496), .Y(n4099) );
   IV110  g608( .A(n4269), .Y(n4939) );
   BF003  g609( .A1(n4308), .A2(n4495), .B1(n4183), .B2(
                           n4494), .Y(n4587) );
   IV110  g610( .A(n4739), .Y(n4737) );
   NO210  g611( .A(n3879), .B(n4143), .Y(n4874) );
   IV110  g612( .A(n4274), .Y(n4937) );
   AN210  g613( .A(A_14_port), .B(B_15_port), .Y(n4872) );
   BF053  g614( .A1(n4327), .A2(n5207), .B1(n4291), .B2(
                           n5174), .Y(n4328) );
   AN210  g615( .A(n4049), .B(n4178), .Y(n4801) );
   IV110  g616( .A(n4278), .Y(n4512) );
   NO210  g617( .A(n3978), .B(n3977), .Y(n4050) );
   NA410  g618( .A(n5007), .B(n4571), .C(n4052), .D(n4053), .Y(
                           n4051) );
   NA210  g619( .A(n4392), .B(n4557), .Y(n5006) );
   NO210  g620( .A(n3976), .B(n4556), .Y(n4573) );
   EX2B0  g621( .A(n5067), .B(n5068), .Y(PRODUCT_16_port) );
   BF003  g622( .A1(n3993), .A2(n4152), .B1(n4714), .B2(
                           n4153), .Y(n5145) );
   EX2B0  g623( .A(n4715), .B(n4151), .Y(n4804) );
   EN2B0  g624( .A(n4716), .B(n4150), .Y(n5153) );
   EN210  g625( .A(n4975), .B(n5190), .Y(n5154) );
   EX2B0  g626( .A(n4149), .B(n5125), .Y(n5105) );
   NA210  g627( .A(n4137), .B(n4139), .Y(n4736) );
   IV110  g628( .A(n4343), .Y(n4341) );
   NO210  g629( .A(n4143), .B(n4142), .Y(n4141) );
   BF053  g630( .A1(n3950), .A2(n3949), .B1(n3882), .B2(
                           n4668), .Y(n4340) );
   NO210  g631( .A(n5062), .B(n4262), .Y(n4140) );
   IV110  g632( .A(n4340), .Y(n4339) );
   NO210  g633( .A(n4140), .B(n4139), .Y(n4138) );
   BF053  g634( .A1(n3880), .A2(n3931), .B1(n3932), .B2(
                           n3944), .Y(n3933) );
   BF053  g635( .A1(n4735), .A2(n4899), .B1(n5132), .B2(
                           n4229), .Y(n4688) );
   IV110  g636( .A(n3933), .Y(n3930) );
   NA210  g637( .A(n4137), .B(n5082), .Y(n5081) );
   NA311  g638( .A(n5065), .B(n4137), .C(n4733), .Y(n4734) );
   NA210  g639( .A(B_3_port), .B(A_10_port), .Y(n3875) );
   NA210  g640( .A(B_1_port), .B(A_13_port), .Y(n3876) );
   NA210  g641( .A(A_8_port), .B(B_6_port), .Y(n3877) );
   IV110  g642( .A(n4691), .Y(n4689) );
   IV110  g643( .A(n4130), .Y(n4131) );
   BF053  g644( .A1(n4466), .A2(n4465), .B1(n4815), .B2(
                           n5021), .Y(n4672) );
   IV110  g645( .A(n4672), .Y(n4671) );
   BF053  g646( .A1(n4669), .A2(n4461), .B1(n4814), .B2(
                           n4594), .Y(n4670) );
   NA210  g647( .A(B_2_port), .B(A_4_port), .Y(n4610) );
   IV110  g648( .A(n4670), .Y(n4668) );
   NO210  g649( .A(n3869), .B(n4187), .Y(n4611) );
   BF053  g650( .A1(n4247), .A2(n4460), .B1(n4812), .B2(
                           n4248), .Y(n4667) );
   NA210  g651( .A(B_2_port), .B(A_6_port), .Y(n4612) );
   IV110  g652( .A(n4667), .Y(n4246) );
   NO210  g653( .A(n3869), .B(n4614), .Y(n4613) );
   BF053  g654( .A1(n4035), .A2(n4032), .B1(n4034), .B2(
                           n4033), .Y(n4245) );
   NA210  g655( .A(B_2_port), .B(A_8_port), .Y(n4615) );
   BF053  g656( .A1(n4463), .A2(n4462), .B1(n4813), .B2(
                           n4590), .Y(n4244) );
   NA210  g657( .A(B_2_port), .B(A_9_port), .Y(n4616) );
   NA210  g658( .A(B_2_port), .B(A_10_port), .Y(n5041) );
   NA210  g659( .A(A_8_port), .B(B_8_port), .Y(n4193) );
   NA210  g660( .A(B_7_port), .B(A_9_port), .Y(n4194) );
   NA210  g661( .A(B_6_port), .B(A_10_port), .Y(n4195) );
   NA210  g662( .A(A_14_port), .B(B_13_port), .Y(n4551) );
   NO210  g663( .A(n4552), .B(n4169), .Y(n4393) );
   NA210  g664( .A(B_13_port), .B(A_15_port), .Y(n4553) );
   NA210  g665( .A(A_14_port), .B(B_14_port), .Y(n4554) );
   NA210  g666( .A(A_13_port), .B(B_15_port), .Y(n4555) );
   NA210  g667( .A(n4176), .B(n4177), .Y(n3977) );
   NA210  g668( .A(n4175), .B(n4393), .Y(n4556) );
   EN210  g669( .A(n4044), .B(n4040), .Y(n4043) );
   IV110  g670( .A(n4725), .Y(n5011) );
   EN210  g671( .A(n4042), .B(n4041), .Y(n4040) );
   EN2B0  g672( .A(n4273), .B(n4643), .Y(n4396) );
   EX2B0  g673( .A(n4039), .B(n4038), .Y(n4037) );
   IV110  g674( .A(n4545), .Y(n4072) );
   EN2B0  g675( .A(n4087), .B(n5075), .Y(n5149) );
   IV110  g676( .A(n4114), .Y(n4502) );
   BF003  g677( .A1(n4938), .A2(n5076), .B1(n4270), .B2(n5073
                           ), .Y(n4095) );
   IV110  g678( .A(n5059), .Y(n4503) );
   BF003  g679( .A1(n4939), .A2(n5074), .B1(n4269), .B2(n4645
                           ), .Y(n5075) );
   NA210  g680( .A(A_4_port), .B(B_13_port), .Y(n4624) );
   EN210  g681( .A(n5040), .B(n4161), .Y(n4096) );
   NA210  g682( .A(A_6_port), .B(B_11_port), .Y(n4625) );
   BF003  g683( .A1(n4940), .A2(n4162), .B1(n3872), .B2(n5077
                           ), .Y(n4161) );
   NA210  g684( .A(B_7_port), .B(A_11_port), .Y(n4626) );
   NA210  g685( .A(B_8_port), .B(A_10_port), .Y(n5051) );
   NA210  g686( .A(B_9_port), .B(A_9_port), .Y(n5052) );
   NA210  g687( .A(A_5_port), .B(B_13_port), .Y(n5053) );
   NA210  g688( .A(A_4_port), .B(B_14_port), .Y(n5054) );
   NA210  g689( .A(B_4_port), .B(A_14_port), .Y(n4629) );
   NA210  g690( .A(B_4_port), .B(A_15_port), .Y(n4630) );
   NA210  g691( .A(n4631), .B(n4792), .Y(n4268) );
   BF003  g692( .A1(n4834), .A2(n4675), .B1(n4280), .B2(
                           n5093), .Y(n4360) );
   EX2B0  g693( .A(n5094), .B(n4281), .Y(n4759) );
   EX210  g694( .A(n4788), .B(n4787), .Y(n4388) );
   EN210  g695( .A(n4791), .B(n4790), .Y(n4789) );
   EX210  g696( .A(n4794), .B(n4793), .Y(n4792) );
   EN2B0  g697( .A(n5215), .B(n4796), .Y(n4795) );
   EN210  g698( .A(n5218), .B(n5217), .Y(n5216) );
   EN2B0  g699( .A(n3860), .B(n3859), .Y(n3858) );
   EX2B0  g700( .A(n3863), .B(n3862), .Y(n3861) );
   BF001  g701( .A1(n4603), .B1(n4602), .B2(n4596), .Y(n4601
                           ) );
   BF003  g702( .A1(n4070), .A2(n4223), .B1(n4547), .B2(
                           n4225), .Y(n4324) );
   NA210  g703( .A(A_2_port), .B(B_6_port), .Y(n4022) );
   BF003  g704( .A1(n4069), .A2(n5169), .B1(n4548), .B2(
                           n5171), .Y(n4738) );
   EN210  g705( .A(n4289), .B(n4738), .Y(n5209) );
   BF003  g706( .A1(n4068), .A2(n5172), .B1(n4290), .B2(
                           n5173), .Y(n5208) );
   IV110  g707( .A(n4058), .Y(n4919) );
   BF053  g708( .A1(n4336), .A2(n4902), .B1(n4621), .B2(
                           n4752), .Y(n4337) );
   IV110  g709( .A(n4065), .Y(n4490) );
   IV110  g710( .A(n4337), .Y(n4335) );
   BF053  g711( .A1(n4203), .A2(n4318), .B1(n3997), .B2(
                           n3969), .Y(n3998) );
   BF053  g712( .A1(n4622), .A2(n4332), .B1(n4623), .B2(
                           n4333), .Y(n4334) );
   BF003  g713( .A1(n4120), .A2(n3998), .B1(n4945), .B2(
                           n5109), .Y(n4552) );
   IV110  g714( .A(n4334), .Y(n4331) );
   NA210  g715( .A(n4556), .B(n3976), .Y(n4053) );
   BF053  g716( .A1(n4624), .A2(n4755), .B1(n4904), .B2(
                           n4903), .Y(n4330) );
   BF053  g717( .A1(n5143), .A2(n3901), .B1(n3973), .B2(
                           n4379), .Y(n3981) );
   NA210  g718( .A(n4989), .B(n3982), .Y(n4987) );
   NA410  g719( .A(n4987), .B(n4603), .C(n4869), .D(n4988), .Y(
                           n4994) );
   IV110  g720( .A(n4544), .Y(n4073) );
   NA210  g721( .A(n4987), .B(n4165), .Y(n4993) );
   EN210  g722( .A(n4901), .B(n4900), .Y(n4899) );
   EN210  g723( .A(n4904), .B(n4903), .Y(n4902) );
   EN210  g724( .A(n4103), .B(n4102), .Y(n4101) );
   EN210  g725( .A(n3955), .B(n3954), .Y(n4905) );
   EN210  g726( .A(n4100), .B(n4099), .Y(n4098) );
   EX210  g727( .A(n3958), .B(n3957), .Y(n3956) );
   EN210  g728( .A(n4097), .B(n4358), .Y(n4357) );
   EN210  g729( .A(n3961), .B(n3960), .Y(n3959) );
   EN210  g730( .A(n4353), .B(n4350), .Y(n4356) );
   EN210  g731( .A(n4355), .B(n4354), .Y(n4353) );
   BF053  g732( .A1(n5139), .A2(n4850), .B1(n4309), .B2(
                           n4487), .Y(n4310) );
   IV110  g733( .A(n4310), .Y(n3903) );
   BF053  g734( .A1(n4912), .A2(n4911), .B1(n5141), .B2(
                           n4856), .Y(n3902) );
   IV110  g735( .A(n3902), .Y(n3901) );
   NA210  g736( .A(n4204), .B(n4380), .Y(n4869) );
   EN210  g737( .A(n4024), .B(n4133), .Y(n4529) );
   BF003  g738( .A1(n4512), .A2(n5080), .B1(n4278), .B2(
                           n5078), .Y(n4127) );
   BF003  g739( .A1(n4511), .A2(n4128), .B1(n4697), .B2(
                           n5079), .Y(n4106) );
   BF003  g740( .A1(n4510), .A2(n4131), .B1(n4700), .B2(
                           n4130), .Y(n4560) );
   BF003  g741( .A1(n4509), .A2(n4561), .B1(n4704), .B2(
                           n4559), .Y(n4531) );
   EX2B0  g742( .A(n4164), .B(n4694), .Y(PRODUCT_24_port) );
   EX210  g743( .A(n4037), .B(n4695), .Y(PRODUCT_13_port) );
   EN2B0  g744( .A(n5081), .B(n4696), .Y(PRODUCT_21_port) );
   EX2B0  g745( .A(n4980), .B(n5105), .Y(PRODUCT_9_port) );
   EN210  g746( .A(n5108), .B(n5107), .Y(n5106) );
   EX210  g747( .A(n5111), .B(n5110), .Y(n5109) );
   EN210  g748( .A(n5114), .B(n5113), .Y(n5112) );
   NO210  g749( .A(n5103), .B(n4705), .Y(n4876) );
   NO210  g750( .A(n3868), .B(n4701), .Y(n4458) );
   NA210  g751( .A(A_2_port), .B(B_8_port), .Y(n4878) );
   BF003  g752( .A1(n4301), .A2(n4586), .B1(n4810), .B2(
                           n4588), .Y(n4468) );
   BF003  g753( .A1(n4300), .A2(n4248), .B1(n4812), .B2(
                           n4589), .Y(n4247) );
   EN210  g754( .A(n4460), .B(n4247), .Y(n4463) );
   BF003  g755( .A1(n4299), .A2(n4590), .B1(n4813), .B2(
                           n4593), .Y(n4462) );
   BF003  g756( .A1(n3893), .A2(n4594), .B1(n4814), .B2(
                           n4595), .Y(n4669) );
   EN210  g757( .A(n4461), .B(n4669), .Y(n4466) );
   BF003  g758( .A1(n3892), .A2(n5021), .B1(n4815), .B2(
                           n5023), .Y(n4465) );
   EN210  g759( .A(n4249), .B(n5214), .Y(n5213) );
   EX210  g760( .A(n4252), .B(n4251), .Y(n4250) );
   EX210  g761( .A(n4255), .B(n4254), .Y(n4253) );
   IV110  g762( .A(n4855), .Y(n4853) );
   IV110  g763( .A(n5063), .Y(n4139) );
   IV110  g764( .A(n5010), .Y(n4210) );
   IV110  g765( .A(n4990), .Y(n4868) );
   IV110  g766( .A(n4991), .Y(n4214) );
   IV110  g767( .A(n4048), .Y(n4641) );
   IV110  g768( .A(n4644), .Y(n5071) );
   BF053  g769( .A1(n5114), .A2(n5113), .B1(n4124), .B2(
                           n4846), .Y(n4842) );
   IV110  g770( .A(n4842), .Y(n4841) );
   BF053  g771( .A1(n4123), .A2(n4839), .B1(n4122), .B2(
                           n4843), .Y(n4840) );
   BF053  g772( .A1(n5088), .A2(n5197), .B1(n4712), .B2(
                           n4757), .Y(n5089) );
   IV110  g773( .A(n5089), .Y(n5087) );
   BF053  g774( .A1(n5199), .A2(n5198), .B1(n4711), .B2(
                           n4346), .Y(n5086) );
   BF003  g775( .A1(n4580), .A2(n4853), .B1(n5140), .B2(
                           n4855), .Y(n4727) );
   IV110  g776( .A(n5086), .Y(n5085) );
   EN210  g777( .A(n4907), .B(n4727), .Y(n4912) );
   BF053  g778( .A1(n5083), .A2(n4776), .B1(n4710), .B2(
                           n4344), .Y(n5084) );
   BF003  g779( .A1(n4579), .A2(n4856), .B1(n5141), .B2(
                           n3904), .Y(n4911) );
   IV110  g780( .A(n5084), .Y(n4666) );
   EN210  g781( .A(n4910), .B(n4729), .Y(n3965) );
   EN210  g782( .A(n5196), .B(n5195), .Y(n4776) );
   BF053  g783( .A1(n4883), .A2(n4882), .B1(n5115), .B2(
                           n4567), .Y(n5001) );
   IV110  g784( .A(n5001), .Y(n5002) );
   EN210  g785( .A(n4470), .B(n5182), .Y(n4475) );
   BF053  g786( .A1(n5005), .A2(n4880), .B1(n4706), .B2(
                           n5004), .Y(n5003) );
   BF003  g787( .A1(n4410), .A2(n4661), .B1(n4193), .B2(
                           n4663), .Y(n4474) );
   IV110  g788( .A(n5003), .Y(n4057) );
   BF003  g789( .A1(n4409), .A2(n4664), .B1(n4194), .B2(
                           n4665), .Y(n4321) );
   BF053  g790( .A1(n4879), .A2(n4878), .B1(n4877), .B2(
                           n4457), .Y(n4058) );
   EN210  g791( .A(n4473), .B(n4321), .Y(n4478) );
   EX2B0  g792( .A(n4177), .B(n4176), .Y(n4175) );
   EN210  g793( .A(n4174), .B(n4173), .Y(n4172) );
   EN210  g794( .A(n4171), .B(n4170), .Y(n4169) );
   EN210  g795( .A(n5200), .B(n5090), .Y(n4976) );
   EN2B0  g796( .A(n4713), .B(n4760), .Y(n5201) );
   EN210  g797( .A(n5197), .B(n5088), .Y(n5202) );
   BF003  g798( .A1(n4417), .A2(n4757), .B1(n4712), .B2(n4758
                           ), .Y(n5088) );
   BF003  g799( .A1(n4418), .A2(n4346), .B1(n4711), .B2(n4348
                           ), .Y(n5198) );
   EN210  g800( .A(n4776), .B(n5083), .Y(n5199) );
   BF003  g801( .A1(n4827), .A2(n4344), .B1(n4710), .B2(n4345
                           ), .Y(n5083) );
   EN210  g802( .A(n4373), .B(n4653), .Y(n4378) );
   EN210  g803( .A(n4376), .B(n4440), .Y(n4779) );
   IV110  g804( .A(n4233), .Y(n4232) );
   BF053  g805( .A1(n4713), .A2(n4760), .B1(n5202), .B2(
                           n5201), .Y(n4231) );
   BF053  g806( .A1(n4283), .A2(n4761), .B1(n5204), .B2(
                           n4976), .Y(n4230) );
   IV110  g807( .A(n4230), .Y(n4229) );
   BF053  g808( .A1(n4475), .A2(n4474), .B1(n4193), .B2(
                           n4661), .Y(n5184) );
   BF053  g809( .A1(n5134), .A2(n4232), .B1(n5182), .B2(
                           n4470), .Y(n5183) );
   BF003  g810( .A1(n4824), .A2(n5158), .B1(n4634), .B2(
                           n5159), .Y(n3862) );
   IV110  g811( .A(n5183), .Y(n5181) );
   IV110  g812( .A(n4699), .Y(n4515) );
   IV110  g813( .A(n4702), .Y(n4517) );
   IV110  g814( .A(n4706), .Y(n4518) );
   IV110  g815( .A(n5119), .Y(n4086) );
   IV110  g816( .A(n4179), .Y(n4080) );
   EX210  g817( .A(n4522), .B(n4519), .Y(PRODUCT_2_port) );
   IV110  g818( .A(n4317), .Y(n4316) );
   EX2B0  g819( .A(n4055), .B(n4054), .Y(PRODUCT_10_port) );
   BF053  g820( .A1(n5136), .A2(n4437), .B1(n4488), .B2(
                           n4906), .Y(n4315) );
   EN210  g821( .A(n4893), .B(n4890), .Y(n3944) );
   IV110  g822( .A(n4315), .Y(n4314) );
   EN210  g823( .A(n4895), .B(n4894), .Y(n4893) );
   BF053  g824( .A1(n5137), .A2(n4847), .B1(n5138), .B2(
                           n4312), .Y(n4313) );
   EN210  g825( .A(n4892), .B(n4891), .Y(n4890) );
   IV110  g826( .A(n4313), .Y(n4311) );
   EX2B0  g827( .A(n4889), .B(n4888), .Y(n4887) );
   EN210  g828( .A(n4886), .B(n4468), .Y(n4467) );
   EN210  g829( .A(n4466), .B(n4465), .Y(n4464) );
   BF053  g830( .A1(n4497), .A2(n3939), .B1(n5121), .B2(
                           n5002), .Y(n4496) );
   EN210  g831( .A(n4463), .B(n4462), .Y(n4461) );
   BF053  g832( .A1(n4893), .A2(n4890), .B1(n4892), .B2(
                           n4891), .Y(n3929) );
   EX2B0  g833( .A(n4298), .B(n4012), .Y(n4010) );
   BF053  g834( .A1(n3881), .A2(n4246), .B1(n3947), .B2(
                           n3946), .Y(n3928) );
   BF003  g835( .A1(n5018), .A2(n4323), .B1(n4717), .B2(
                           n4325), .Y(n4854) );
   BF053  g836( .A1(n3878), .A2(n4243), .B1(n3926), .B2(
                           n3945), .Y(n3927) );
   NA210  g837( .A(A_5_port), .B(B_9_port), .Y(n3878) );
   BF003  g838( .A1(n5017), .A2(n4326), .B1(n4718), .B2(
                           n4328), .Y(n4851) );
   NA210  g839( .A(A_2_port), .B(B_12_port), .Y(n4891) );
   IV110  g840( .A(n3927), .Y(n3925) );
   NA210  g841( .A(n4459), .B(n4036), .Y(n4892) );
   BF003  g842( .A1(n5016), .A2(n4737), .B1(n4719), .B2(
                           n4739), .Y(n4848) );
   NO210  g843( .A(n5103), .B(n3879), .Y(n4895) );
   BF053  g844( .A1(n4282), .A2(n5096), .B1(n4364), .B2(
                           n4363), .Y(n3924) );
   NO210  g845( .A(n3868), .B(n4811), .Y(n4894) );
   EN210  g846( .A(n4720), .B(n4848), .Y(n4685) );
   NA210  g847( .A(A_3_port), .B(B_11_port), .Y(n3880) );
   NA210  g848( .A(A_4_port), .B(B_10_port), .Y(n3881) );
   NA210  g849( .A(A_5_port), .B(B_14_port), .Y(n4111) );
   NA210  g850( .A(A_4_port), .B(B_15_port), .Y(n4112) );
   NA210  g851( .A(A_6_port), .B(B_13_port), .Y(n4113) );
   IV110  g852( .A(n4244), .Y(n4243) );
   BF053  g853( .A1(n4816), .A2(n5024), .B1(n4241), .B2(
                           n4464), .Y(n4242) );
   EX2B0  g854( .A(n4867), .B(n4395), .Y(PRODUCT_25_port) );
   EX210  g855( .A(n4525), .B(n4396), .Y(PRODUCT_3_port) );
   BF003  g856( .A1(n4397), .A2(n4602), .B1(n4167), .B2(
                           n4398), .Y(PRODUCT_22_port) );
   NA210  g857( .A(B_5_port), .B(A_11_port), .Y(n4196) );
   EX210  g858( .A(n4799), .B(n4798), .Y(n4797) );
   NA210  g859( .A(B_4_port), .B(A_12_port), .Y(n4197) );
   EX2B0  g860( .A(n4797), .B(n4801), .Y(n4800) );
   NA210  g861( .A(B_2_port), .B(A_14_port), .Y(n4198) );
   EX2B0  g862( .A(n4983), .B(n4802), .Y(PRODUCT_11_port) );
   NA210  g863( .A(B_7_port), .B(A_10_port), .Y(n4617) );
   EN2B0  g864( .A(n4569), .B(n4803), .Y(PRODUCT_29_port) );
   NO210  g865( .A(n4698), .B(n5048), .Y(n4618) );
   EX2B0  g866( .A(n4977), .B(n4804), .Y(PRODUCT_7_port) );
   NA210  g867( .A(A_8_port), .B(B_9_port), .Y(n4619) );
   NA210  g868( .A(A_7_port), .B(B_10_port), .Y(n4620) );
   NA210  g869( .A(A_14_port), .B(B_10_port), .Y(n4203) );
   NO210  g870( .A(n3964), .B(n3965), .Y(n4382) );
   NA210  g871( .A(n4913), .B(n4384), .Y(n4204) );
   EX2B0  g872( .A(n4874), .B(n4875), .Y(n4873) );
   NA210  g873( .A(n4895), .B(n4894), .Y(n4768) );
   EX210  g874( .A(n4872), .B(n4873), .Y(n4799) );
   NA210  g875( .A(A_3_port), .B(B_12_port), .Y(n4288) );
   EX210  g876( .A(n4141), .B(n4642), .Y(n4638) );
   NA210  g877( .A(A_4_port), .B(B_11_port), .Y(n4707) );
   IV110  g878( .A(n4688), .Y(n4690) );
   NA210  g879( .A(A_7_port), .B(B_8_port), .Y(n4708) );
   IV110  g880( .A(n4914), .Y(n3964) );
   NA210  g881( .A(A_8_port), .B(B_7_port), .Y(n4709) );
   EX210  g882( .A(n4985), .B(n4984), .Y(n4983) );
   EX2B0  g883( .A(n4982), .B(n4981), .Y(n4980) );
   EX2B0  g884( .A(n4979), .B(n4978), .Y(n4977) );
   BF053  g885( .A1(n4531), .A2(n4532), .B1(n4704), .B2(
                           n4561), .Y(n4996) );
   EX210  g886( .A(n4976), .B(n5204), .Y(n5203) );
   IV110  g887( .A(n4996), .Y(n4997) );
   EX210  g888( .A(n5202), .B(n5201), .Y(n5200) );
   BF053  g889( .A1(n4999), .A2(n4881), .B1(n5116), .B2(
                           n4563), .Y(n4998) );
   BF001  g890( .A1(n4048), .B1(n4052), .B2(n4806), .Y(n3867
                           ) );
   EN210  g891( .A(n5199), .B(n5198), .Y(n5197) );
   BF051  g892( .A1(n5065), .B1(n4210), .B2(n4732), .Y(n3866
                           ) );
   IV110  g893( .A(n4998), .Y(n5000) );
   NA311  g894( .A(n4573), .B(n4941), .C(n4639), .Y(n4803) );
   IV110  g895( .A(n4280), .Y(n4834) );
   IV110  g896( .A(n5041), .Y(n4302) );
   IV110  g897( .A(n5102), .Y(n5100) );
   NA210  g898( .A(A_8_port), .B(B_15_port), .Y(n5138) );
   IV110  g899( .A(n4610), .Y(n4304) );
   OR210  g900( .A(n4795), .B(n4268), .Y(n4632) );
   NA210  g901( .A(A_9_port), .B(B_14_port), .Y(n5137) );
   NO210  g902( .A(n5216), .B(n4632), .Y(n4603) );
   IV110  g903( .A(n4810), .Y(n4301) );
   NA210  g904( .A(B_3_port), .B(A_14_port), .Y(n4633) );
   NA210  g905( .A(B_3_port), .B(A_15_port), .Y(n4634) );
   NA210  g906( .A(n4261), .B(n4260), .Y(n4264) );
   NO210  g907( .A(n4263), .B(n4264), .Y(n4635) );
   NA210  g908( .A(B_2_port), .B(A_15_port), .Y(n4636) );
   NA210  g909( .A(n4641), .B(n4052), .Y(n4805) );
   NA210  g910( .A(n4797), .B(n4801), .Y(n4637) );
   NA210  g911( .A(n4995), .B(n4987), .Y(n4395) );
   EN2B0  g912( .A(n4261), .B(n4260), .Y(n4259) );
   NO210  g913( .A(n5006), .B(n4574), .Y(n4600) );
   EX210  g914( .A(n4264), .B(n4263), .Y(n4262) );
   BF006  g915( .A1(n4598), .A2(n4599), .B1(n4571), .B2(
                           n4573), .Y(n4597) );
   EX210  g916( .A(n4266), .B(n4259), .Y(n4265) );
   BF003  g917( .A1(n4873), .A2(n4872), .B1(n4875), .B2(
                           n4874), .Y(n4871) );
   BF006  g918( .A1(n4870), .A2(n4165), .B1(n4869), .B2(
                           n4868), .Y(n4867) );
   NA210  g919( .A(n4596), .B(n4168), .Y(n4167) );
   NO210  g920( .A(n4166), .B(n4165), .Y(n4164) );
   NO210  g921( .A(n5104), .B(n5103), .Y(PRODUCT_0_port) );
   IV110  g922( .A(n4330), .Y(n4329) );
   EN210  g923( .A(n5106), .B(n4425), .Y(n5111) );
   BF053  g924( .A1(n3921), .A2(n4905), .B1(n4620), .B2(
                           n3922), .Y(n3923) );
   BF003  g925( .A1(n4405), .A2(n4001), .B1(n4119), .B2(
                           n4002), .Y(n5110) );
   IV110  g926( .A(n3923), .Y(n3920) );
   IV110  g927( .A(n4543), .Y(n4074) );
   EX2B0  g928( .A(n4120), .B(n3998), .Y(n4945) );
   NA310  g929( .A(n4869), .B(n4868), .C(n4987), .Y(n4992) );
   BF053  g930( .A1(n3918), .A2(n4370), .B1(n5051), .B2(
                           n4751), .Y(n3919) );
   IV110  g931( .A(n4541), .Y(n4075) );
   BF003  g932( .A1(n4404), .A2(n3999), .B1(n4121), .B2(
                           n4000), .Y(n4170) );
   BF051  g933( .A1(n4214), .B1(n4986), .B2(n4398), .Y(n4806
                           ) );
   BF053  g934( .A1(n4371), .A2(n4372), .B1(n5052), .B2(
                           n4748), .Y(n3917) );
   IV110  g935( .A(n4540), .Y(n4076) );
   BF003  g936( .A1(n4403), .A2(n4843), .B1(n4122), .B2(
                           n4845), .Y(n4839) );
   NA210  g937( .A(n4047), .B(n4389), .Y(n4052) );
   IV110  g938( .A(n4546), .Y(n4071) );
   IV110  g939( .A(n4547), .Y(n4070) );
   IV110  g940( .A(n4292), .Y(n5020) );
   IV110  g941( .A(n4291), .Y(n4067) );
   EN210  g942( .A(n4352), .B(n4351), .Y(n4350) );
   IV110  g943( .A(n4593), .Y(n4590) );
   EN210  g944( .A(n4349), .B(n3943), .Y(n3942) );
   BF053  g945( .A1(n4353), .A2(n4350), .B1(n4352), .B2(
                           n4351), .Y(n4589) );
   EN210  g946( .A(n3941), .B(n3940), .Y(n3939) );
   BF003  g947( .A1(n4820), .A2(n4311), .B1(n4199), .B2(
                           n4313), .Y(n3898) );
   BF053  g948( .A1(n4183), .A2(n4495), .B1(n4587), .B2(
                           n4098), .Y(n4588) );
   EN210  g949( .A(n4200), .B(n3898), .Y(n3968) );
   EN210  g950( .A(n3935), .B(n4884), .Y(n3938) );
   IV110  g951( .A(n4328), .Y(n4326) );
   IV110  g952( .A(n4588), .Y(n4586) );
   BF053  g953( .A1(n4547), .A2(n4223), .B1(n4324), .B2(
                           n5210), .Y(n4325) );
   EN210  g954( .A(n3937), .B(n3936), .Y(n3935) );
   IV110  g955( .A(n4325), .Y(n4323) );
   BF053  g956( .A1(n4161), .A2(n5040), .B1(n3872), .B2(
                           n4162), .Y(n4163) );
   BF053  g957( .A1(n4321), .A2(n4473), .B1(n4194), .B2(
                           n4664), .Y(n4322) );
   IV110  g958( .A(n4322), .Y(n4320) );
   BF053  g959( .A1(n4254), .A2(n4255), .B1(n4617), .B2(
                           n4320), .Y(n4319) );
   IV110  g960( .A(n4607), .Y(n4307) );
   IV110  g961( .A(n4319), .Y(n3913) );
   BF003  g962( .A1(n4086), .A2(n4919), .B1(n5119), .B2(
                           n4058), .Y(n4920) );
   EN210  g963( .A(n3938), .B(n4920), .Y(n3941) );
   BF003  g964( .A1(n4085), .A2(n4057), .B1(n5120), .B2(
                           n5003), .Y(n3940) );
   BF003  g965( .A1(n4084), .A2(n5002), .B1(n5121), .B2(
                           n5001), .Y(n4497) );
   EN210  g966( .A(n3939), .B(n4497), .Y(n4349) );
   NA210  g967( .A(A_12_port), .B(B_9_port), .Y(n4293) );
   NO210  g968( .A(n4277), .B(n4807), .Y(n4294) );
   NA210  g969( .A(A_12_port), .B(B_6_port), .Y(n4295) );
   NO210  g970( .A(n4285), .B(n4277), .Y(n4296) );
   NA210  g971( .A(A_14_port), .B(B_6_port), .Y(n4297) );
   NA210  g972( .A(n4449), .B(n4026), .Y(n4879) );
   NA210  g973( .A(A_3_port), .B(B_7_port), .Y(n4706) );
   NA210  g974( .A(A_4_port), .B(B_6_port), .Y(n5115) );
   NA210  g975( .A(B_5_port), .B(A_5_port), .Y(n5116) );
   NA210  g976( .A(B_4_port), .B(A_7_port), .Y(n5117) );
   NA210  g977( .A(n4876), .B(n4458), .Y(n3934) );
   NA210  g978( .A(A_2_port), .B(B_9_port), .Y(n4885) );
   NO210  g979( .A(n5103), .B(n4142), .Y(n4367) );
   NO210  g980( .A(n3868), .B(n3879), .Y(n4366) );
   NA210  g981( .A(A_2_port), .B(B_13_port), .Y(n4767) );
   EN210  g982( .A(n4258), .B(n4257), .Y(n4256) );
   EX210  g983( .A(n4679), .B(n4678), .Y(n4677) );
   EN210  g984( .A(n4682), .B(n4681), .Y(n4680) );
   EN210  g985( .A(n4685), .B(n4684), .Y(n4683) );
   EN210  g986( .A(n4023), .B(n4022), .Y(n4021) );
   EN210  g987( .A(n4480), .B(n4479), .Y(n4686) );
   EN210  g988( .A(n4020), .B(n4019), .Y(n4018) );
   EN210  g989( .A(n4483), .B(n4482), .Y(n4481) );
   EN210  g990( .A(n4017), .B(n4965), .Y(n4964) );
   EN210  g991( .A(n4486), .B(n4485), .Y(n4484) );
   IV110  g992( .A(n4840), .Y(n4838) );
   BF053  g993( .A1(n4428), .A2(n3966), .B1(n5144), .B2(
                           n3903), .Y(n4837) );
   IV110  g994( .A(n4837), .Y(n4427) );
   IV110  g995( .A(n4625), .Y(n3987) );
   BF053  g996( .A1(n4425), .A2(n5106), .B1(n4118), .B2(
                           n4427), .Y(n4426) );
   IV110  g997( .A(n4624), .Y(n3988) );
   IV110  g998( .A(n4426), .Y(n4424) );
   IV110  g999( .A(n4754), .Y(n4332) );
   BF053  g1000( .A1(n4125), .A2(n4424), .B1(n4422), .B2(
                           n5112), .Y(n4423) );
   IV110  g1001( .A(n4621), .Y(n3990) );
   BF053  g1002( .A1(n5196), .A2(n5195), .B1(n4709), .B2(
                           n4341), .Y(n4665) );
   EN210  g1003( .A(n4484), .B(n5142), .Y(n5218) );
   EN210  g1004( .A(n4253), .B(n4429), .Y(n4788) );
   BF003  g1005( .A1(n4578), .A2(n4007), .B1(n4205), .B2(
                           n4009), .Y(n4787) );
   BF003  g1006( .A1(n4577), .A2(n4954), .B1(n4206), .B2(
                           n4955), .Y(n4790) );
   EN210  g1007( .A(n4256), .B(n4015), .Y(n4791) );
   EN210  g1008( .A(n4677), .B(n4013), .Y(n4387) );
   IV110  g1009( .A(n4222), .Y(n4221) );
   BF053  g1010( .A1(n4219), .A2(n4780), .B1(n4543), .B2(
                           n4652), .Y(n4220) );
   IV110  g1011( .A(n4220), .Y(n5174) );
   BF053  g1012( .A1(n5037), .A2(n5034), .B1(n5039), .B2(
                           n5038), .Y(n4059) );
   BF003  g1013( .A1(n3996), .A2(n4666), .B1(n4195), .B2(
                           n5084), .Y(n4477) );
   BF003  g1014( .A1(n3995), .A2(n5085), .B1(n4196), .B2(
                           n5086), .Y(n4008) );
   EN210  g1015( .A(n4476), .B(n4008), .Y(n4898) );
   BF003  g1016( .A1(n3994), .A2(n5087), .B1(n4197), .B2(
                           n5089), .Y(n4897) );
   EN210  g1017( .A(n4896), .B(n5160), .Y(n4901) );
   EN210  g1018( .A(n4198), .B(n5091), .Y(n4900) );
   BF053  g1019( .A1(n3876), .A2(n4762), .B1(n4763), .B2(
                           n4362), .Y(n4764) );
   IV110  g1020( .A(n4764), .Y(n4761) );
   BF003  g1021( .A1(n4281), .A2(n5094), .B1(n4759), .B2(
                           n4359), .Y(n4760) );
   EN210  g1022( .A(n4789), .B(n5164), .Y(n3863) );
   BF053  g1023( .A1(n4472), .A2(n4471), .B1(n4192), .B2(
                           n4660), .Y(n5180) );
   EX2B0  g1024( .A(n4385), .B(n5162), .Y(n4260) );
   BF053  g1025( .A1(n5178), .A2(n4045), .B1(n4189), .B2(
                           n4234), .Y(n5179) );
   BF003  g1026( .A1(n4823), .A2(n5156), .B1(n4636), .B2(
                           n5157), .Y(n5155) );
   IV110  g1027( .A(n5179), .Y(n5177) );
   EX2B0  g1028( .A(n3861), .B(n5061), .Y(n4693) );
   EN210  g1029( .A(n3858), .B(n5155), .Y(n4691) );
   BF003  g1030( .A1(n4822), .A2(n3901), .B1(n5143), .B2(
                           n3902), .Y(n3973) );
   BF003  g1031( .A1(n4821), .A2(n3903), .B1(n5144), .B2(
                           n4310), .Y(n4428) );
   IV110  g1032( .A(n4496), .Y(n4498) );
   EN210  g1033( .A(n4035), .B(n4032), .Y(n4460) );
   BF053  g1034( .A1(n3941), .A2(n3940), .B1(n5120), .B2(
                           n4057), .Y(n4916) );
   EN210  g1035( .A(n4459), .B(n4036), .Y(n4035) );
   IV110  g1036( .A(n4916), .Y(n4917) );
   EN210  g1037( .A(n4034), .B(n4033), .Y(n4032) );
   BF053  g1038( .A1(n4920), .A2(n3938), .B1(n5119), .B2(
                           n4919), .Y(n4918) );
   IV110  g1039( .A(n4918), .Y(n4921) );
   EN210  g1040( .A(n5126), .B(n4148), .Y(n4055) );
   BF053  g1041( .A1(n4885), .A2(n3934), .B1(n3935), .B2(
                           n4884), .Y(n4922) );
   BF003  g1042( .A1(n5015), .A2(n4740), .B1(n4721), .B2(
                           n4741), .Y(n4684) );
   EN210  g1043( .A(n4683), .B(n4851), .Y(n4480) );
   BF003  g1044( .A1(n4742), .A2(n5014), .B1(n4743), .B2(
                           n4722), .Y(n4479) );
   EN210  g1045( .A(n4686), .B(n4854), .Y(n4483) );
   BF003  g1046( .A1(n4744), .A2(n5013), .B1(n4745), .B2(
                           n4723), .Y(n4482) );
   NA210  g1047( .A(A_13_port), .B(B_7_port), .Y(n4114) );
   IV110  g1048( .A(n4857), .Y(n4448) );
   NA210  g1049( .A(A_12_port), .B(B_8_port), .Y(n4115) );
   BF053  g1050( .A1(n4445), .A2(n4777), .B1(n5060), .B2(
                           n4446), .Y(n4447) );
   NA210  g1051( .A(B_9_port), .B(A_11_port), .Y(n4116) );
   IV110  g1052( .A(n4447), .Y(n4444) );
   NA210  g1053( .A(B_10_port), .B(A_10_port), .Y(n4539) );
   BF053  g1054( .A1(n4778), .A2(n4779), .B1(n4107), .B2(
                           n3916), .Y(n4443) );
   NA210  g1055( .A(A_7_port), .B(B_13_port), .Y(n4540) );
   IV110  g1056( .A(n4443), .Y(n4442) );
   NA210  g1057( .A(A_6_port), .B(B_14_port), .Y(n4541) );
   NA210  g1058( .A(A_5_port), .B(B_15_port), .Y(n4542) );
   NA210  g1059( .A(A_11_port), .B(B_14_port), .Y(n5070) );
   NA210  g1060( .A(A_10_port), .B(B_15_port), .Y(n4117) );
   NA210  g1061( .A(A_13_port), .B(B_12_port), .Y(n4118) );
   EN210  g1062( .A(n4806), .B(n4805), .Y(PRODUCT_26_port) );
   EX210  g1063( .A(n5203), .B(n3864), .Y(PRODUCT_15_port) );
   NO210  g1064( .A(n3868), .B(n5118), .Y(n4354) );
   NA210  g1065( .A(A_3_port), .B(B_9_port), .Y(n4179) );
   NA210  g1066( .A(A_4_port), .B(B_8_port), .Y(n4180) );
   IV110  g1067( .A(n4711), .Y(n4418) );
   NA210  g1068( .A(A_5_port), .B(B_7_port), .Y(n4181) );
   NA210  g1069( .A(B_5_port), .B(A_12_port), .Y(n4205) );
   NA210  g1070( .A(A_6_port), .B(B_6_port), .Y(n4182) );
   IV110  g1071( .A(n4710), .Y(n4827) );
   NA210  g1072( .A(B_5_port), .B(A_7_port), .Y(n4183) );
   NA210  g1073( .A(B_5_port), .B(A_13_port), .Y(n4206) );
   AN210  g1074( .A(A_3_port), .B(B_3_port), .Y(n4184) );
   IV110  g1075( .A(n4709), .Y(n4828) );
   NA210  g1076( .A(B_3_port), .B(A_4_port), .Y(n4185) );
   NA210  g1077( .A(B_5_port), .B(A_14_port), .Y(n4207) );
   IV110  g1078( .A(n4708), .Y(n4829) );
   NA210  g1079( .A(B_5_port), .B(A_15_port), .Y(n4208) );
   IV110  g1080( .A(n4707), .Y(n4830) );
   NA210  g1081( .A(n4796), .B(n5215), .Y(n5217) );
   IV110  g1082( .A(n4602), .Y(n4398) );
   NA210  g1083( .A(B_6_port), .B(A_9_port), .Y(n4710) );
   IV110  g1084( .A(n4209), .Y(n4211) );
   NA210  g1085( .A(B_5_port), .B(A_10_port), .Y(n4711) );
   IV110  g1086( .A(A_9_port), .Y(n5048) );
   IV110  g1087( .A(A_7_port), .Y(n4614) );
   IV110  g1088( .A(A_5_port), .Y(n4187) );
   BF053  g1089( .A1(n4206), .A2(n4954), .B1(n4791), .B2(
                           n4790), .Y(n4953) );
   IV110  g1090( .A(n4953), .Y(n4952) );
   BF053  g1091( .A1(n4207), .A2(n4952), .B1(n4386), .B2(
                           n4387), .Y(n4951) );
   NA210  g1092( .A(A_10_port), .B(B_13_port), .Y(n5136) );
   IV110  g1093( .A(n4589), .Y(n4248) );
   NA210  g1094( .A(A_12_port), .B(B_11_port), .Y(n5135) );
   IV110  g1095( .A(n4813), .Y(n4299) );
   NA210  g1096( .A(B_8_port), .B(A_15_port), .Y(n4726) );
   IV110  g1097( .A(n4814), .Y(n3893) );
   NA210  g1098( .A(B_7_port), .B(A_15_port), .Y(n4725) );
   IV110  g1099( .A(n4815), .Y(n3892) );
   IV110  g1100( .A(n5069), .Y(n4408) );
   NA210  g1101( .A(A_14_port), .B(B_8_port), .Y(n4724) );
   NA210  g1102( .A(n4990), .B(n4988), .Y(n3865) );
   IV110  g1103( .A(n4816), .Y(n3891) );
   IV110  g1104( .A(n4124), .Y(n4402) );
   OR210  g1105( .A(n3982), .B(n4989), .Y(n4995) );
   IV110  g1106( .A(n4122), .Y(n4403) );
   NA210  g1107( .A(n4798), .B(n4799), .Y(n4642) );
   IV110  g1108( .A(n4551), .Y(n3986) );
   BF003  g1109( .A1(n4520), .A2(n4521), .B1(n4522), .B2(
                           n4519), .Y(n4643) );
   IV110  g1110( .A(n4549), .Y(n4399) );
   BF053  g1111( .A1(n4273), .A2(n4643), .B1(n4396), .B2(
                           n4525), .Y(n4644) );
   BF001  g1112( .A1(n5010), .B1(n5009), .B2(n5008), .Y(
                           PRODUCT_18_port) );
   NA210  g1113( .A(n4956), .B(n4528), .Y(n4023) );
   NA210  g1114( .A(n5007), .B(n5006), .Y(n4575) );
   NA210  g1115( .A(A_3_port), .B(B_5_port), .Y(n4699) );
   NA210  g1116( .A(B_4_port), .B(A_5_port), .Y(n4700) );
   BF003  g1117( .A1(n4067), .A2(n5174), .B1(n4291), .B2(
                           n4220), .Y(n4327) );
   NO210  g1118( .A(n5103), .B(n4701), .Y(n4449) );
   EN210  g1119( .A(n5207), .B(n4327), .Y(n5212) );
   NO210  g1120( .A(n3868), .B(n4698), .Y(n4026) );
   BF003  g1121( .A1(n5020), .A2(n4221), .B1(n4292), .B2(
                           n4222), .Y(n5211) );
   EN210  g1122( .A(n4123), .B(n4839), .Y(n5114) );
   BF003  g1123( .A1(n4402), .A2(n4846), .B1(n4124), .B2(
                           n3894), .Y(n5113) );
   BF003  g1124( .A1(n4401), .A2(n4424), .B1(n4125), .B2(
                           n4426), .Y(n4422) );
   EN210  g1125( .A(n5112), .B(n4422), .Y(n4171) );
   BF003  g1126( .A1(n4400), .A2(n4421), .B1(n4126), .B2(
                           n4423), .Y(n4420) );
   IV110  g1127( .A(n4290), .Y(n4068) );
   BF053  g1128( .A1(n4718), .A2(n4326), .B1(n4851), .B2(
                           n4683), .Y(n4852) );
   IV110  g1129( .A(n4548), .Y(n4069) );
   IV110  g1130( .A(n4852), .Y(n4850) );
   BF003  g1131( .A1(n4303), .A2(n5100), .B1(n4616), .B2(
                           n5102), .Y(n5099) );
   BF053  g1132( .A1(n4719), .A2(n4737), .B1(n4720), .B2(
                           n4848), .Y(n4849) );
   BF003  g1133( .A1(n4302), .A2(n5098), .B1(n5041), .B2(
                           n5101), .Y(n4970) );
   IV110  g1134( .A(n4849), .Y(n4847) );
   EN210  g1135( .A(n4533), .B(n4157), .Y(n4979) );
   BF053  g1136( .A1(n4721), .A2(n4740), .B1(n4685), .B2(
                           n4684), .Y(n4438) );
   EX2B0  g1137( .A(n4239), .B(n5042), .Y(n5193) );
   EN2B0  g1138( .A(n5044), .B(n5194), .Y(n4978) );
   EX2B0  g1139( .A(n5045), .B(n5192), .Y(n5190) );
   EN2B0  g1140( .A(n4536), .B(n4154), .Y(n4982) );
   EN2B0  g1141( .A(n5046), .B(n5191), .Y(n4981) );
   IV110  g1142( .A(n4163), .Y(n4160) );
   EN210  g1143( .A(n5055), .B(n4862), .Y(n3961) );
   BF053  g1144( .A1(n4610), .A2(n4160), .B1(n4973), .B2(
                           n4974), .Y(n4159) );
   BF003  g1145( .A1(n4932), .A2(n4335), .B1(n5056), .B2(
                           n4337), .Y(n4859) );
   BF003  g1146( .A1(n4611), .A2(n4159), .B1(n4157), .B2(
                           n4533), .Y(n4158) );
   IV110  g1147( .A(n4616), .Y(n4303) );
   EN210  g1148( .A(n3959), .B(n4859), .Y(n4369) );
   BF053  g1149( .A1(n4257), .A2(n4258), .B1(n4626), .B2(
                           n3913), .Y(n3912) );
   BF053  g1150( .A1(n4027), .A2(n4028), .B1(n4612), .B2(
                           n4158), .Y(n4156) );
   IV110  g1151( .A(n4812), .Y(n4300) );
   BF003  g1152( .A1(n4931), .A2(n4338), .B1(n5057), .B2(
                           n4747), .Y(n3963) );
   IV110  g1153( .A(n3912), .Y(n3911) );
   BF003  g1154( .A1(n4154), .A2(n4536), .B1(n4613), .B2(
                           n4156), .Y(n4155) );
   IV110  g1155( .A(n3876), .Y(n4833) );
   BF003  g1156( .A1(n4930), .A2(n3920), .B1(n5058), .B2(
                           n3923), .Y(n3914) );
   BF053  g1157( .A1(n5059), .A2(n3911), .B1(n4678), .B2(
                           n4679), .Y(n3910) );
   IV110  g1158( .A(n3880), .Y(n3886) );
   IV110  g1159( .A(n4288), .Y(n4831) );
   IV110  g1160( .A(n4190), .Y(n4412) );
   IV110  g1161( .A(n4620), .Y(n3991) );
   NO210  g1162( .A(n4277), .B(n4143), .Y(n4298) );
   NA210  g1163( .A(A_12_port), .B(B_10_port), .Y(n4717) );
   NA210  g1164( .A(B_12_port), .B(A_10_port), .Y(n4718) );
   NA210  g1165( .A(A_8_port), .B(B_14_port), .Y(n4719) );
   NA210  g1166( .A(A_7_port), .B(B_15_port), .Y(n4720) );
   NA210  g1167( .A(n3981), .B(n3980), .Y(n4390) );
   NO210  g1168( .A(n4391), .B(n4390), .Y(n4557) );
   NA210  g1169( .A(n4558), .B(n3972), .Y(n3983) );
   NA410  g1170( .A(n4869), .B(n4987), .C(n4596), .D(n4988), 
                           .Y(n4986) );
   NA210  g1171( .A(n4381), .B(n4382), .Y(n4989) );
   NA210  g1172( .A(A_4_port), .B(B_9_port), .Y(n4813) );
   NA210  g1173( .A(A_5_port), .B(B_8_port), .Y(n4814) );
   NA210  g1174( .A(A_6_port), .B(B_7_port), .Y(n4815) );
   NA210  g1175( .A(A_7_port), .B(B_6_port), .Y(n4816) );
   NA210  g1176( .A(B_4_port), .B(A_9_port), .Y(n3874) );
   NA210  g1177( .A(A_3_port), .B(B_15_port), .Y(n5055) );
   NA210  g1178( .A(A_6_port), .B(B_12_port), .Y(n5056) );
   NA210  g1179( .A(A_7_port), .B(B_11_port), .Y(n5057) );
   NA210  g1180( .A(A_8_port), .B(B_10_port), .Y(n5058) );
   NA210  g1181( .A(A_12_port), .B(B_7_port), .Y(n5059) );
   EN210  g1182( .A(n4963), .B(n4962), .Y(n4961) );
   EN210  g1183( .A(n4527), .B(n4957), .Y(n4960) );
   EN210  g1184( .A(n4959), .B(n4958), .Y(n4957) );
   EN210  g1185( .A(n4956), .B(n4528), .Y(n4527) );
   EX2B0  g1186( .A(n4094), .B(n4526), .Y(PRODUCT_5_port) );
   EN210  g1187( .A(n4091), .B(n4088), .Y(n4525) );
   NA210  g1188( .A(A_0_port), .B(B_1_port), .Y(n4271) );
   EX2B0  g1189( .A(n4524), .B(n4523), .Y(n4522) );
   NA210  g1190( .A(A_1_port), .B(B_0_port), .Y(n4272) );
   NO210  g1191( .A(n4271), .B(n4272), .Y(n4521) );
   IV110  g1192( .A(n4423), .Y(n4421) );
   IV110  g1193( .A(n5052), .Y(n4935) );
   IV110  g1194( .A(n5057), .Y(n4931) );
   IV110  g1195( .A(n5056), .Y(n4932) );
   IV110  g1196( .A(n5054), .Y(n4933) );
   IV110  g1197( .A(n5053), .Y(n4934) );
   IV110  g1198( .A(n5058), .Y(n4930) );
   EN210  g1199( .A(n4098), .B(n4587), .Y(n4103) );
   EN210  g1200( .A(n4454), .B(n4560), .Y(n4538) );
   EX210  g1201( .A(n4184), .B(n4059), .Y(n4061) );
   BF053  g1202( .A1(n4540), .A2(n4647), .B1(n4781), .B2(
                           n4782), .Y(n5173) );
   IV110  g1203( .A(n5173), .Y(n5172) );
   BF053  g1204( .A1(n4542), .A2(n5170), .B1(n4541), .B2(
                           n4649), .Y(n5171) );
   IV110  g1205( .A(B_11_port), .Y(n5118) );
   IV110  g1206( .A(n5171), .Y(n5169) );
   IV110  g1207( .A(B_3_port), .Y(n3870) );
   BF053  g1208( .A1(n5205), .A2(n5206), .B1(n4116), .B2(
                           n4442), .Y(n5168) );
   IV110  g1209( .A(B_12_port), .Y(n5124) );
   IV110  g1210( .A(n5168), .Y(n5167) );
   IV110  g1211( .A(B_14_port), .Y(n3879) );
   BF053  g1212( .A1(n4361), .A2(n4360), .B1(n4280), .B2(
                           n4675), .Y(n4758) );
   IV110  g1213( .A(n4758), .Y(n4757) );
   BF053  g1214( .A1(n4347), .A2(n3951), .B1(n4279), .B2(
                           n4673), .Y(n4348) );
   IV110  g1215( .A(n4348), .Y(n4346) );
   BF053  g1216( .A1(n3952), .A2(n3953), .B1(n3877), .B2(
                           n4240), .Y(n4345) );
   IV110  g1217( .A(n4345), .Y(n4344) );
   BF053  g1218( .A1(n3883), .A2(n4671), .B1(n4342), .B2(
                           n3948), .Y(n4343) );
   IV110  g1219( .A(n3917), .Y(n3916) );
   BF053  g1220( .A1(n5058), .A2(n3920), .B1(n3914), .B2(
                           n3962), .Y(n3915) );
   IV110  g1221( .A(n3915), .Y(n4866) );
   EN210  g1222( .A(n4906), .B(n4488), .Y(n4487) );
   EN210  g1223( .A(n4909), .B(n4908), .Y(n4907) );
   EN210  g1224( .A(n4912), .B(n4911), .Y(n4910) );
   BF003  g1225( .A1(n4915), .A2(n4914), .B1(n3965), .B2(
                           n3964), .Y(n4913) );
   EN210  g1226( .A(n3968), .B(n3967), .Y(n3966) );
   EX2B0  g1227( .A(n5127), .B(n4147), .Y(n4802) );
   BF053  g1228( .A1(n5117), .A2(n4997), .B1(n4924), .B2(
                           n3942), .Y(n4923) );
   EN210  g1229( .A(n5128), .B(n4146), .Y(n5152) );
   IV110  g1230( .A(n4923), .Y(n4925) );
   EX210  g1231( .A(n5129), .B(n4145), .Y(n4695) );
   BF053  g1232( .A1(n5029), .A2(n4101), .B1(n4609), .B2(
                           n4493), .Y(n5030) );
   EN210  g1233( .A(n5130), .B(n4144), .Y(n5147) );
   EX210  g1234( .A(n5131), .B(n5092), .Y(n3864) );
   BF003  g1235( .A1(n3992), .A2(n5181), .B1(n4619), .B2(
                           n5183), .Y(n3957) );
   BF003  g1236( .A1(n3991), .A2(n3922), .B1(n4620), .B2(
                           n5180), .Y(n3921) );
   BF053  g1237( .A1(n4440), .A2(n4376), .B1(n4108), .B2(
                           n4866), .Y(n4441) );
   IV110  g1238( .A(n4441), .Y(n4439) );
   BF053  g1239( .A1(n4109), .A2(n4448), .B1(n4377), .B2(
                           n4378), .Y(n4656) );
   IV110  g1240( .A(n4656), .Y(n4655) );
   BF053  g1241( .A1(n4110), .A2(n4858), .B1(n4653), .B2(
                           n4373), .Y(n4654) );
   NA210  g1242( .A(A_14_port), .B(B_11_port), .Y(n4119) );
   NA210  g1243( .A(A_2_port), .B(B_11_port), .Y(n4033) );
   NO210  g1244( .A(n4705), .B(n4143), .Y(n4120) );
   NA210  g1245( .A(n4355), .B(n4354), .Y(n4034) );
   NA210  g1246( .A(B_11_port), .B(A_15_port), .Y(n4121) );
   NO210  g1247( .A(n5103), .B(n4811), .Y(n4459) );
   NA210  g1248( .A(A_12_port), .B(B_14_port), .Y(n4122) );
   NO210  g1249( .A(n3868), .B(n5124), .Y(n4036) );
   NA210  g1250( .A(A_11_port), .B(B_15_port), .Y(n4123) );
   NA210  g1251( .A(A_3_port), .B(B_10_port), .Y(n4812) );
   NA210  g1252( .A(A_13_port), .B(B_13_port), .Y(n4124) );
   NA210  g1253( .A(A_14_port), .B(B_12_port), .Y(n4125) );
   BF053  g1254( .A1(n4699), .A2(n4134), .B1(n4133), .B2(
                           n4024), .Y(n4132) );
   IV110  g1255( .A(n4132), .Y(n4135) );
   BF053  g1256( .A1(n4021), .A2(n4018), .B1(n4023), .B2(
                           n4022), .Y(n4136) );
   NO210  g1257( .A(n3870), .B(n4187), .Y(n4186) );
   NA210  g1258( .A(B_3_port), .B(A_6_port), .Y(n4188) );
   NA210  g1259( .A(B_0_port), .B(A_14_port), .Y(n5130) );
   NO210  g1260( .A(n5104), .B(n4143), .Y(n5131) );
   NA210  g1261( .A(B_1_port), .B(A_15_port), .Y(n5132) );
   IV110  g1262( .A(n3929), .Y(n4238) );
   NO210  g1263( .A(n3870), .B(n4285), .Y(n5133) );
   NO210  g1264( .A(n5218), .B(n5217), .Y(n4627) );
   NA210  g1265( .A(A_7_port), .B(B_9_port), .Y(n5134) );
   IV110  g1266( .A(n4286), .Y(n4832) );
   NA210  g1267( .A(A_5_port), .B(B_11_port), .Y(n4189) );
   NO210  g1268( .A(n3871), .B(n4285), .Y(n4628) );
   NA210  g1269( .A(A_1_port), .B(B_15_port), .Y(n4044) );
   IV110  g1270( .A(n4714), .Y(n3993) );
   NA210  g1271( .A(A_3_port), .B(B_13_port), .Y(n4190) );
   IV110  g1272( .A(n4197), .Y(n3994) );
   IV110  g1273( .A(n4196), .Y(n3995) );
   BF056  g1274( .A1(n4215), .A2(n4570), .B1(n4051), .B2(
                           n4214), .Y(n4598) );
   BF052  g1275( .A1(n4217), .B1(n4574), .B2(n5006), .B3(
                           n4216), .Y(n4599) );
   EX210  g1276( .A(n4638), .B(n4637), .Y(n4218) );
   IV110  g1277( .A(n4951), .Y(n4950) );
   BF053  g1278( .A1(n4794), .A2(n4793), .B1(n4208), .B2(
                           n4950), .Y(n4796) );
   NO210  g1279( .A(n4627), .B(n4383), .Y(n4212) );
   IV110  g1280( .A(n4608), .Y(n4306) );
   BF053  g1281( .A1(n4197), .A2(n5087), .B1(n4898), .B2(
                           n4897), .Y(n4949) );
   IV110  g1282( .A(n4609), .Y(n4305) );
   BF003  g1283( .A1(n4947), .A2(n4388), .B1(n4628), .B2(
                           n4949), .Y(n4948) );
   IV110  g1284( .A(n4183), .Y(n4308) );
   BF053  g1285( .A1(n4629), .A2(n4948), .B1(n5164), .B2(
                           n4789), .Y(n4946) );
   IV110  g1286( .A(n4182), .Y(n4077) );
   BF003  g1287( .A1(n4499), .A2(n4439), .B1(n4539), .B2(
                           n4441), .Y(n4224) );
   NO210  g1288( .A(n3868), .B(n4277), .Y(n4528) );
   BF003  g1289( .A1(n4076), .A2(n4647), .B1(n4540), .B2(
                           n4648), .Y(n4781) );
   NO210  g1290( .A(n3868), .B(n3873), .Y(n4965) );
   BF003  g1291( .A1(n4075), .A2(n4649), .B1(n4541), .B2(
                           n4651), .Y(n5170) );
   EN210  g1292( .A(n4542), .B(n5170), .Y(n4782) );
   BF003  g1293( .A1(n4074), .A2(n4652), .B1(n4543), .B2(
                           n4654), .Y(n4219) );
   BF053  g1294( .A1(n4190), .A2(n4756), .B1(n5175), .B2(
                           n4043), .Y(n5176) );
   IV110  g1295( .A(n5176), .Y(n4755) );
   BF051  g1296( .A1(n4042), .B1(n4044), .B2(n4040), .Y(n4754
                           ) );
   NA210  g1297( .A(A_13_port), .B(B_9_port), .Y(n4723) );
   NA210  g1298( .A(B_11_port), .B(A_11_port), .Y(n4722) );
   NA210  g1299( .A(A_9_port), .B(B_13_port), .Y(n4721) );
   IV110  g1300( .A(A_15_port), .Y(n4143) );
   IV110  g1301( .A(B_2_port), .Y(n3869) );
   IV110  g1302( .A(A_0_port), .Y(n5103) );
   NO210  g1303( .A(n5104), .B(n4285), .Y(n5129) );
   IV110  g1304( .A(A_1_port), .Y(n3868) );
   IV110  g1305( .A(n4118), .Y(n4406) );
   NA210  g1306( .A(B_0_port), .B(A_12_port), .Y(n5128) );
   BF053  g1307( .A1(n4091), .A2(n4088), .B1(n4090), .B2(
                           n4089), .Y(n4645) );
   IV110  g1308( .A(B_0_port), .Y(n5104) );
   IV110  g1309( .A(n4125), .Y(n4401) );
   BF053  g1310( .A1(n5150), .A2(n5149), .B1(n4274), .B2(
                           n5071), .Y(n4646) );
   IV110  g1311( .A(n4126), .Y(n4400) );
   IV110  g1312( .A(n4554), .Y(n3984) );
   IV110  g1313( .A(n4553), .Y(n3985) );
   BF003  g1314( .A1(n4829), .A2(n4339), .B1(n4708), .B2(
                           n4340), .Y(n4662) );
   EN210  g1315( .A(n4773), .B(n4662), .Y(n5196) );
   BF003  g1316( .A1(n4828), .A2(n4341), .B1(n4709), .B2(
                           n4343), .Y(n5195) );
   NA210  g1317( .A(A_2_port), .B(B_7_port), .Y(n4451) );
   EN210  g1318( .A(n5210), .B(n4324), .Y(n4249) );
   NA210  g1319( .A(n4020), .B(n4019), .Y(n4452) );
   BF003  g1320( .A1(n5019), .A2(n5167), .B1(n4293), .B2(
                           n5168), .Y(n5214) );
   NA210  g1321( .A(A_3_port), .B(B_6_port), .Y(n4702) );
   EN210  g1322( .A(n5213), .B(n5165), .Y(n4252) );
   NA210  g1323( .A(B_5_port), .B(A_4_port), .Y(n4703) );
   EX2B0  g1324( .A(n4294), .B(n4431), .Y(n4429) );
   NA210  g1325( .A(B_4_port), .B(A_6_port), .Y(n4704) );
   EN2B0  g1326( .A(n4295), .B(n4430), .Y(n4015) );
   IV110  g1327( .A(n4438), .Y(n4437) );
   IV110  g1328( .A(n4645), .Y(n5074) );
   BF053  g1329( .A1(n4722), .A2(n4742), .B1(n4480), .B2(
                           n4479), .Y(n4436) );
   IV110  g1330( .A(n4275), .Y(n4936) );
   IV110  g1331( .A(n4436), .Y(n4435) );
   EX2B0  g1332( .A(n5047), .B(n5189), .Y(n5187) );
   IV110  g1333( .A(n4270), .Y(n4938) );
   EN210  g1334( .A(n4966), .B(n5099), .Y(n4985) );
   BF053  g1335( .A1(n4433), .A2(n4481), .B1(n4724), .B2(
                           n4746), .Y(n4434) );
   EN210  g1336( .A(n4369), .B(n3963), .Y(n3962) );
   IV110  g1337( .A(n5077), .Y(n4162) );
   EN210  g1338( .A(n4372), .B(n4371), .Y(n4370) );
   IV110  g1339( .A(n4434), .Y(n4432) );
   EN210  g1340( .A(n4375), .B(n4374), .Y(n4373) );
   IV110  g1341( .A(n5078), .Y(n5080) );
   EN210  g1342( .A(n4378), .B(n4377), .Y(n4376) );
   EN210  g1343( .A(n4779), .B(n4778), .Y(n4777) );
   EN210  g1344( .A(n4782), .B(n4781), .Y(n4780) );
   EN210  g1345( .A(n4785), .B(n4784), .Y(n4783) );
   EN210  g1346( .A(n3934), .B(n4885), .Y(n4884) );
   EN210  g1347( .A(n3962), .B(n3914), .Y(n4372) );
   EN210  g1348( .A(n4370), .B(n3918), .Y(n4258) );
   EN210  g1349( .A(n3956), .B(n4750), .Y(n4255) );
   BF003  g1350( .A1(n4929), .A2(n4320), .B1(n4617), .B2(
                           n4322), .Y(n4254) );
   BF003  g1351( .A1(n4928), .A2(n3913), .B1(n4626), .B2(
                           n4319), .Y(n4257) );
   IV110  g1352( .A(n4622), .Y(n3989) );
   IV110  g1353( .A(n4665), .Y(n4664) );
   IV110  g1354( .A(n5060), .Y(n4927) );
   BF053  g1355( .A1(n4708), .A2(n4339), .B1(n4662), .B2(
                           n4773), .Y(n4663) );
   NA310  g1356( .A(n4733), .B(n5010), .C(n4640), .Y(n3900) );
   IV110  g1357( .A(n4663), .Y(n4661) );
   BF056  g1358( .A1(n5063), .A2(n3900), .B1(n5065), .B2(
                           n4140), .Y(n4696) );
   BF003  g1359( .A1(n4287), .A2(n3928), .B1(n4659), .B2(
                           n4770), .Y(n4660) );
   BF053  g1360( .A1(n4199), .A2(n4311), .B1(n4200), .B2(
                           n3898), .Y(n3899) );
   BF053  g1361( .A1(n4288), .A2(n4238), .B1(n4657), .B2(
                           n4769), .Y(n4658) );
   IV110  g1362( .A(n3899), .Y(n3897) );
   BF053  g1363( .A1(n4201), .A2(n4314), .B1(n3968), .B2(
                           n3967), .Y(n3896) );
   IV110  g1364( .A(n3896), .Y(n3895) );
   IV110  g1365( .A(n4195), .Y(n3996) );
   BF053  g1366( .A1(n5107), .A2(n5108), .B1(n5069), .B2(
                           n3895), .Y(n3894) );
   NO210  g1367( .A(n4380), .B(n4204), .Y(n4165) );
   NA210  g1368( .A(n4383), .B(n4627), .Y(n4990) );
   NA410  g1369( .A(n4993), .B(n4992), .C(n4994), .D(n4995), 
                           .Y(n4991) );
   OR210  g1370( .A(n3979), .B(n3983), .Y(n4047) );
   NO210  g1371( .A(n4389), .B(n4047), .Y(n4048) );
   EN210  g1372( .A(n4481), .B(n4433), .Y(n4486) );
   EN210  g1373( .A(n4775), .B(n4774), .Y(n4773) );
   BF003  g1374( .A1(n4802), .A2(n4983), .B1(n5127), .B2(
                           n4147), .Y(n4146) );
   EX210  g1375( .A(n4772), .B(n4771), .Y(n4770) );
   BF003  g1376( .A1(n5011), .A2(n3905), .B1(n4725), .B2(
                           n3906), .Y(n4485) );
   EN210  g1377( .A(n4365), .B(n4368), .Y(n4769) );
   BF053  g1378( .A1(n5152), .A2(n5151), .B1(n5128), .B2(
                           n4146), .Y(n4145) );
   EN210  g1379( .A(n4768), .B(n4767), .Y(n4368) );
   BF003  g1380( .A1(n4585), .A2(n4432), .B1(n4726), .B2(
                           n4434), .Y(n4729) );
   EN210  g1381( .A(n4367), .B(n4366), .Y(n4365) );
   BF003  g1382( .A1(n4695), .A2(n4037), .B1(n5129), .B2(
                           n4145), .Y(n4144) );
   BF003  g1383( .A1(n4584), .A2(n4435), .B1(n5135), .B2(
                           n4436), .Y(n4908) );
   BF003  g1384( .A1(n4437), .A2(n4583), .B1(n4438), .B2(
                           n5136), .Y(n4488) );
   BF003  g1385( .A1(n4582), .A2(n4847), .B1(n5137), .B2(
                           n4849), .Y(n4312) );
   EN210  g1386( .A(n5138), .B(n4312), .Y(n4906) );
   NA210  g1387( .A(B_8_port), .B(A_11_port), .Y(n5060) );
   NA210  g1388( .A(B_9_port), .B(A_10_port), .Y(n4107) );
   NA210  g1389( .A(B_10_port), .B(A_9_port), .Y(n4108) );
   NA210  g1390( .A(A_8_port), .B(B_11_port), .Y(n4109) );
   NA210  g1391( .A(A_7_port), .B(B_12_port), .Y(n4110) );
   NA210  g1392( .A(n5061), .B(n3861), .Y(n4266) );
   NO210  g1393( .A(n4259), .B(n4266), .Y(n5062) );
   NA210  g1394( .A(n4262), .B(n5062), .Y(n5063) );
   NO210  g1395( .A(n4690), .B(n4691), .Y(n4692) );
   AN210  g1396( .A(n4693), .B(n4692), .Y(n5064) );

endmodule

module csa_mult_n17_m17_1

       ( A_16_port, A_15_port, A_14_port, A_13_port, A_12_port, A_11_port, 
         A_10_port, A_9_port, A_8_port, A_7_port, A_6_port, A_5_port, A_4_port,
         A_3_port, A_2_port, A_1_port, A_0_port, B_16_port, B_15_port, 
         B_14_port, B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, 
         B_8_port, B_7_port, B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, 
         B_1_port, B_0_port, CTL, PRODUCT_33_port, 
         PRODUCT_32_port, PRODUCT_31_port, PRODUCT_30_port, PRODUCT_29_port, 
         PRODUCT_28_port, PRODUCT_27_port, PRODUCT_26_port, PRODUCT_25_port, 
         PRODUCT_24_port, PRODUCT_23_port, PRODUCT_22_port, PRODUCT_21_port, 
         PRODUCT_20_port, PRODUCT_19_port, PRODUCT_18_port, PRODUCT_17_port, 
         PRODUCT_16_port, PRODUCT_15_port, PRODUCT_14_port, PRODUCT_13_port, 
         PRODUCT_12_port, PRODUCT_11_port, PRODUCT_10_port, PRODUCT_9_port, 
         PRODUCT_8_port, PRODUCT_7_port, PRODUCT_6_port, PRODUCT_5_port, 
         PRODUCT_4_port, PRODUCT_3_port, PRODUCT_2_port, PRODUCT_1_port, 
         PRODUCT_0_port);
 
input    A_16_port, A_15_port, A_14_port, A_13_port, A_12_port, A_11_port,
         A_10_port, A_9_port, A_8_port, A_7_port, A_6_port, A_5_port, A_4_port,
         A_3_port, A_2_port, A_1_port, A_0_port, B_16_port, B_15_port,
         B_14_port, B_13_port, B_12_port, B_11_port, B_10_port, B_9_port,
         B_8_port, B_7_port, B_6_port, B_5_port, B_4_port, B_3_port, B_2_port,
         B_1_port, B_0_port, CTL;

output   PRODUCT_33_port,
         PRODUCT_32_port, PRODUCT_31_port, PRODUCT_30_port, PRODUCT_29_port,
         PRODUCT_28_port, PRODUCT_27_port, PRODUCT_26_port, PRODUCT_25_port,
         PRODUCT_24_port, PRODUCT_23_port, PRODUCT_22_port, PRODUCT_21_port,
         PRODUCT_20_port, PRODUCT_19_port, PRODUCT_18_port, PRODUCT_17_port,
         PRODUCT_16_port, PRODUCT_15_port, PRODUCT_14_port, PRODUCT_13_port,
         PRODUCT_12_port, PRODUCT_11_port, PRODUCT_10_port, PRODUCT_9_port,
         PRODUCT_8_port, PRODUCT_7_port, PRODUCT_6_port, PRODUCT_5_port,
         PRODUCT_4_port, PRODUCT_3_port, PRODUCT_2_port, PRODUCT_1_port,
         PRODUCT_0_port;
  
wire  n5709, n5708, n5707, n5706, n5705, n5704, n5703, n5702, n5701, 
      n5700, n5629, n5628, n5627, n5626, n5625, n5624, n5623, n5622, n5621, 
      n5620, n5549, n5548, n5547, n5546, n5545, n5544, n5543, n5542, n5541, 
      n5540, n5469, n5468, n5467, n6519, n5466, n6518, n5465, n6517, n5464, 
      n6516, n5463, n6515, n5462, n6514, n5461, n6513, n5460, n6512, n6511, 
      n6510, n5389, n5388, n5387, n6439, n5386, n6438, n5385, n6437, n5384, 
      n6436, n5383, n6435, n5382, n6434, n5381, n6433, n5380, n6432, n6431, 
      n6430, n6359, n6358, n6357, n6356, n6355, n6354, n6353, n6352, n6351, 
      n6350, n6279, n6278, n6277, n6276, n6275, n6274, n6273, n6272, n6271, 
      n6270, n6199, n6198, n6197, n6196, n6195, n6194, n6193, n6192, n6191, 
      n6190, n5819, n5818, n5817, n5816, n5815, n5814, n5813, n5812, n5811, 
      n5810, n5739, n5738, n5737, n5736, n5735, n5734, n5733, n5732, n5731, 
      n5730, n5659, n5658, n5657, n5656, n5655, n5654, n5653, n5652, n5651, 
      n5650, n5579, n5578, n5577, n5576, n5575, n5574, n5573, n5572, n5571, 
      n5570, n5499, n5498, n5497, n6549, n5496, n6548, n5495, n6547, n5494, 
      n6546, n5493, n6545, n5492, n6544, n5491, n6543, n5490, n6542, n6541, 
      n6540, n6469, n6468, n6467, n6466, n6465, n6464, n6463, n6462, n6461, 
      n6460, n6389, n6388, n6387, n6386, n6385, n6384, n6383, n6382, n6381, 
      n6380, n5929, n5928, n5927, n5926, n5925, n5924, n5923, n5922, n5921, 
      n5920, n5849, n5848, n5847, n5846, n5845, n5844, n5843, n5842, n5841, 
      n5840, n5769, n5768, n5767, n5766, n5765, n5764, n5763, n5762, n5761, 
      n5760, n5689, n5688, n5687, n5686, n5685, n5684, n5683, n5682, n5681, 
      n5680, n6579, n6578, n6577, n6576, n6575, n6574, n6573, n6572, n6571, 
      n6570, n6499, n6498, n6497, n6496, n6495, n6494, n6493, n6492, n6491, 
      n6490, n6019, n6018, n6017, n6016, n6015, n6014, n6013, n6012, n6011, 
      n6010, n5959, n5958, n5957, n5956, n5955, n5954, n5953, n5952, n5951, 
      n5950, n5879, n5878, n5877, n5876, n5875, n5874, n5873, n5872, n5871, 
      n5870, n5799, n5798, n5797, n5796, n5795, n5794, n5793, n5792, n5791, 
      n5790, n5319, n5318, n5317, n5316, n5315, n5314, n5313, n5312, n5311, 
      n5310, n5239, n5238, n5237, n5236, n5235, n5234, n5233, n5232, n5231, 
      n5230, n6209, n6208, n6207, n6206, n6205, n6204, n6203, n6202, n6201, 
      n6200, n6129, n6128, n6127, n6126, n6125, n6124, n6123, n6122, n6121, 
      n6120, n6049, n6048, n6047, n6046, n6045, n6044, n6043, n6042, n6041, 
      n6040, n5989, n5988, n5987, n5986, n5985, n5984, n5983, n5982, n5981, 
      n5980, n5509, n5508, n5507, n5506, n5505, n5504, n5503, n5502, n5501, 
      n5500, n5429, n5428, n5427, n5426, n5425, n5424, n5423, n5422, n5421, 
      n5420, n5349, n5348, n5347, n5346, n5345, n5344, n5343, n5342, n5341, 
      n5340, n5269, n5268, n5267, n6319, n5266, n6318, n5265, n6317, n5264, 
      n6316, n5263, n6315, n5262, n6314, n5261, n6313, n5260, n6312, n6311, 
      n6310, n6239, n6238, n6237, n6236, n6235, n6234, n6233, n6232, n6231, 
      n6230, n6159, n6158, n6157, n6156, n6155, n6154, n6153, n6152, n6151, 
      n6150, n6079, n6078, n6077, n6076, n6075, n6074, n6073, n6072, n6071, 
      n6070, n5619, n5618, n5617, n5616, n5615, n5614, n5613, n5612, n5611, 
      n5610, n5539, n5538, n5537, n5536, n5535, n5534, n5533, n5532, n5531, 
      n5530, n5459, n5458, n5457, n6509, n5456, n6508, n5455, n6507, n5454, 
      n6506, n5453, n6505, n5452, n6504, n5451, n6503, n5450, n6502, n6501, 
      n6500, n5379, n5378, n5377, n6429, n5376, n6428, n5375, n6427, n5374, 
      n6426, n5373, n6425, n5372, n6424, n5371, n6423, n5370, n6422, n6421, 
      n6420, n5299, n5298, n5297, n6349, n5296, n6348, n5295, n6347, n5294, 
      n6346, n5293, n6345, n5292, n6344, n5291, n6343, n5290, n6342, n6341, 
      n6340, n6269, n6268, n6267, n6266, n6265, n6264, n6263, n6262, n6261, 
      n6260, n6189, n6188, n6187, n6186, n6185, n6184, n6183, n6182, n6181, 
      n6180, n5809, n5808, n5807, n5806, n5805, n5804, n5803, n5802, n5801, 
      n5800, n5729, n5728, n5727, n5726, n5725, n5724, n5723, n5722, n5721, 
      n5720, n5649, n5648, n5647, n5646, n5645, n5644, n5643, n5642, n5641, 
      n5640, n5569, n5568, n5567, n5566, n5565, n5564, n5563, n5562, n5561, 
      n5560, n5489, n5488, n5487, n6539, n5486, n6538, n5485, n6537, n5484, 
      n6536, n5483, n6535, n5482, n6534, n5481, n6533, n5480, n6532, n6531, 
      n6530, n6459, n6458, n6457, n6456, n6455, n6454, n6453, n6452, n6451, 
      n6450, n6379, n6378, n6377, n6376, n6375, n6374, n6373, n6372, n6371, 
      n6370, n6299, n6298, n6297, n6296, n6295, n6294, n6293, n6292, n6291, 
      n6290, n5919, n5918, n5917, n5916, n5915, n5914, n5913, n5912, n5911, 
      n5910, n5839, n5838, n5837, n5836, n5835, n5834, n5833, n5832, n5831, 
      n5830, n5759, n5758, n5757, n5756, n5755, n5754, n5753, n5752, n5751, 
      n5750, n5679, n5678, n5677, n5676, n5675, n5674, n5673, n5672, n5671, 
      n5670, n5599, n5598, n5597, n5596, n5595, n5594, n5593, n5592, n5591, 
      n5590, n6569, n6568, n6567, n6566, n6565, n6564, n6563, n6562, n6561, 
      n6560, n6489, n6488, n6487, n6486, n6485, n6484, n6483, n6482, n6481, 
      n6480, n6009, n6008, n6007, n6006, n6005, n6004, n6003, n6002, n6001, 
      n6000, n5949, n5948, n5947, n5946, n5945, n5944, n5943, n5942, n5941, 
      n5940, n5869, n5868, n5867, n5866, n5865, n5864, n5863, n5862, n5861, 
      n5860, n5789, n5788, n5787, n5786, n5785, n5784, n5783, n5782, n5781, 
      n5780, n5309, n5308, n5307, n5306, n5305, n5304, n5303, n5302, n5301, 
      n5300, n5229, n5228, n5227, n5226, n5225, n5224, n5223, n5222, n5221, 
      n5220, n6592, n6591, n6590, n6119, n6118, n6117, n6116, n6115, n6114, 
      n6113, n6112, n6111, n6110, n6039, n6038, n6037, n6036, n6035, n6034, 
      n6033, n6032, n6031, n6030, n5979, n5978, n5977, n5976, n5975, n5974, 
      n5973, n5972, n5971, n5970, n5899, n5898, n5897, n5896, n5895, n5894, 
      n5893, n5892, n5891, n5890, n5419, n5418, n5417, n5416, n5415, n5414, 
      n5413, n5412, n5411, n5410, n5339, n5338, n5337, n5336, n5335, n5334, 
      n5333, n5332, n5331, n5330, n5259, n5258, n5257, n6309, n5256, n6308, 
      n5255, n6307, n5254, n6306, n5253, n6305, n5252, n6304, n5251, n6303, 
      n5250, n6302, n6301, n6300, n6229, n6228, n6227, n6226, n6225, n6224, 
      n6223, n6222, n6221, n6220, n6149, n6148, n6147, n6146, n6145, n6144, 
      n6143, n6142, n6141, n6140, n6069, n6068, n6067, n6066, n6065, n6064, 
      n6063, n6062, n6061, n6060, n5609, n5608, n5607, n5606, n5605, n5604, 
      n5603, n5602, n5601, n5600, n5529, n5528, n5527, n5526, n5525, n5524, 
      n5523, n5522, n5521, n5520, n5449, n5448, n5447, n5446, n5445, n5444, 
      n5443, n5442, n5441, n5440, n5369, n5368, n5367, n6419, n5366, n6418, 
      n5365, n6417, n5364, n6416, n5363, n6415, n5362, n6414, n5361, n6413, 
      n5360, n6412, n6411, n6410, n5289, n5288, n5287, n6339, n5286, n6338, 
      n5285, n6337, n5284, n6336, n5283, n6335, n5282, n6334, n5281, n6333, 
      n5280, n6332, n6331, n6330, n6259, n6258, n6257, n6256, n6255, n6254, 
      n6253, n6252, n6251, n6250, n6179, n6178, n6177, n6176, n6175, n6174, 
      n6173, n6172, n6171, n6170, n6099, n6098, n6097, n6096, n6095, n6094, 
      n6093, n6092, n6091, n6090, n5719, n5718, n5717, n5716, n5715, n5714, 
      n5713, n5712, n5711, n5710, n5639, n5638, n5637, n5636, n5635, n5634, 
      n5633, n5632, n5631, n5630, n5559, n5558, n5557, n5556, n5555, n5554, 
      n5553, n5552, n5551, n5550, n5479, n5478, n5477, n6529, n5476, n6528, 
      n5475, n6527, n5474, n6526, n5473, n6525, n5472, n6524, n5471, n6523, 
      n5470, n6522, n6521, n6520, n5399, n5398, n5397, n6449, n5396, n6448, 
      n5395, n6447, n5394, n6446, n5393, n6445, n5392, n6444, n5391, n6443, 
      n5390, n6442, n6441, n6440, n6369, n6368, n6367, n6366, n6365, n6364, 
      n6363, n6362, n6361, n6360, n6289, n6288, n6287, n6286, n6285, n6284, 
      n6283, n6282, n6281, n6280, n5909, n5908, n5907, n5906, n5905, n5904, 
      n5903, n5902, n5901, n5900, n5829, n5828, n5827, n5826, n5825, n5824, 
      n5823, n5822, n5821, n5820, n5749, n5748, n5747, n5746, n5745, n5744, 
      n5743, n5742, n5741, n5740, n5669, n5668, n5667, n5666, n5665, n5664, 
      n5663, n5662, n5661, n5660, n5589, n5588, n5587, n5586, n5585, n5584, 
      n5583, n5582, n5581, n5580, n6559, n6558, n6557, n6556, n6555, n6554, 
      n6553, n6552, n6551, n6550, n6479, n6478, n6477, n6476, n6475, n6474, 
      n6473, n6472, n6471, n6470, n6399, n6398, n6397, n6396, n6395, n6394, 
      n6393, n6392, n6391, n6390, n5939, n5938, n5937, n5936, n5935, n5934, 
      n5933, n5932, n5931, n5930, n5859, n5858, n5857, n5856, n5855, n5854, 
      n5853, n5852, n5851, n5850, n5779, n5778, n5777, n5776, n5775, n5774, 
      n5773, n5772, n5771, n5770, n5699, n5698, n5697, n5696, n5695, n5694, 
      n5693, n5692, n5691, n5690, n5219, n6589, n6588, n6587, n6586, n6585, 
      n6584, n6583, n6582, n6581, n6580, n6109, n6108, n6107, n6106, n6105, 
      n6104, n6103, n6102, n6101, n6100, n6029, n6028, n6027, n6026, n6025, 
      n6024, n6023, n6022, n6021, n6020, n5969, n5968, n5967, n5966, n5965, 
      n5964, n5963, n5962, n5961, n5960, n5889, n5888, n5887, n5886, n5885, 
      n5884, n5883, n5882, n5881, n5880, n5409, n5408, n5407, n5406, n5405, 
      n5404, n5403, n5402, n5401, n5400, n5329, n5328, n5327, n5326, n5325, 
      n5324, n5323, n5322, n5321, n5320, n5249, n5248, n5247, n5246, n5245, 
      n5244, n5243, n5242, n5241, n5240, n6219, n6218, n6217, n6216, n6215, 
      n6214, n6213, n6212, n6211, n6210, n6139, n6138, n6137, n6136, n6135, 
      n6134, n6133, n6132, n6131, n6130, n6059, n6058, n6057, n6056, n6055, 
      n6054, n6053, n6052, n6051, n6050, n5999, n5998, n5997, n5996, n5995, 
      n5994, n5993, n5992, n5991, n5990, n5519, n5518, n5517, n5516, n5515, 
      n5514, n5513, n5512, n5511, n5510, n5439, n5438, n5437, n5436, n5435, 
      n5434, n5433, n5432, n5431, n5430, n5359, n5358, n5357, n6409, n5356, 
      n6408, n5355, n6407, n5354, n6406, n5353, n6405, n5352, n6404, n5351, 
      n6403, n5350, n6402, n6401, n6400, n5279, n5278, n5277, n6329, n5276, 
      n6328, n5275, n6327, n5274, n6326, n5273, n6325, n5272, n6324, n5271, 
      n6323, n5270, n6322, n6321, n6320, n6249, n6248, n6247, n6246, n6245, 
      n6244, n6243, n6242, n6241, n6240, n6169, n6168, n6167, n6166, n6165, 
      n6164, n6163, n6162, n6161, n6160, n6089, n6088, n6087, n6086, n6085, 
      n6084, n6083, n6082, n6081, n6080;

   NA210  g1( .A(A_15_port), .B(B_8_port), .Y(n6093) );
   NO210  g2( .A(n6094), .B(n6052), .Y(n5329) );
   NA210  g3( .A(A_10_port), .B(B_14_port), .Y(n6095) );
   IV110  g4( .A(n6036), .Y(n5718) );
   NA210  g5( .A(A_9_port), .B(B_15_port), .Y(n6509) );
   IV110  g6( .A(n5981), .Y(n5452) );
   NA210  g7( .A(A_11_port), .B(B_13_port), .Y(n6510) );
   IV110  g8( .A(n6416), .Y(n5360) );
   NA210  g9( .A(B_12_port), .B(A_12_port), .Y(n6511) );
   IV110  g10( .A(n6568), .Y(n5711) );
   NA210  g11( .A(A_4_port), .B(B_5_port), .Y(n5647) );
   EN210  g12( .A(n5621), .B(n5805), .Y(n5626) );
   AN210  g13( .A(A_3_port), .B(B_3_port), .Y(n5648) );
   EN210  g14( .A(n5741), .B(n5598), .Y(n6583) );
   NA210  g15( .A(A_4_port), .B(B_3_port), .Y(n5649) );
   EN210  g16( .A(n5317), .B(n5817), .Y(n6580) );
   NO210  g17( .A(n5644), .B(n6173), .Y(n6066) );
   BF003  g18( .A1(n5955), .A2(n5701), .B1(n5569), .B2(
                           n5703), .Y(n6153) );
   EN210  g19( .A(n6267), .B(n5282), .Y(n6154) );
   BF003  g20( .A1(n5954), .A2(n5284), .B1(n5986), .B2(
                           n5700), .Y(n6579) );
   EN210  g21( .A(n5322), .B(n5321), .Y(n5320) );
   EN210  g22( .A(n5740), .B(n5324), .Y(n5323) );
   EX210  g23( .A(n5743), .B(n5742), .Y(n5741) );
   EN210  g24( .A(n5746), .B(n5745), .Y(n5744) );
   EN210  g25( .A(n5749), .B(n5748), .Y(n5747) );
   EN210  g26( .A(n6148), .B(n6147), .Y(n6146) );
   EN210  g27( .A(n6151), .B(n6150), .Y(n6149) );
   EN210  g28( .A(n6249), .B(n6248), .Y(n6247) );
   EX210  g29( .A(n6154), .B(n6153), .Y(n6152) );
   EN210  g30( .A(n6246), .B(n6245), .Y(n6244) );
   NA210  g31( .A(n6003), .B(n5224), .Y(n6011) );
   NO210  g32( .A(n6001), .B(n5221), .Y(n5507) );
   OR210  g33( .A(n5579), .B(n6161), .Y(n5510) );
   NA410  g34( .A(n5510), .B(n6385), .C(n5258), .D(n6011), 
                           .Y(n5259) );
   NA210  g35( .A(n5510), .B(n5506), .Y(n5257) );
   NA310  g36( .A(n5258), .B(n6004), .C(n5510), .Y(n5256) );
   IV110  g37( .A(n6081), .Y(n5251) );
   NA410  g38( .A(n5257), .B(n5256), .C(n5259), .D(n5509), 
                           .Y(n6240) );
   IV110  g39( .A(n6080), .Y(n5252) );
   NA311  g40( .A(n5580), .B(n5533), .C(n6240), .Y(n5255) );
   BF003  g41( .A1(n5948), .A2(n6216), .B1(n5664), .B2(
                           n6217), .Y(n5628) );
   BF053  g42( .A1(n5839), .A2(n6254), .B1(n5838), .B2(
                           n5835), .Y(n5513) );
   BF003  g43( .A1(n5947), .A2(n6218), .B1(n5665), .B2(
                           n6220), .Y(n5378) );
   BF053  g44( .A1(n6185), .A2(n6466), .B1(n5511), .B2(
                           n6255), .Y(n5512) );
   EN210  g45( .A(n5627), .B(n5378), .Y(n6048) );
   BF003  g46( .A1(n5946), .A2(n6221), .B1(n5666), .B2(
                           n6222), .Y(n6047) );
   BF003  g47( .A1(n6195), .A2(n6223), .B1(n5667), .B2(
                           n6225), .Y(n5383) );
   EN210  g48( .A(n6046), .B(n5383), .Y(n6051) );
   BF003  g49( .A1(n6194), .A2(n5265), .B1(n5668), .B2(
                           n5266), .Y(n6050) );
   EN210  g50( .A(n6049), .B(n5801), .Y(n6054) );
   EX2B0  g51( .A(n6524), .B(n6523), .Y(PRODUCT_8_port) );
   EN210  g52( .A(n6525), .B(n6385), .Y(PRODUCT_19_port) );
   BF002  g53( .A1(n5538), .B1(n5928), .B2(n5926), .B3(
                           n6526), .Y(n6362) );
   BF001  g54( .A1(n5944), .B1(n5415), .B2(n5941), .Y(
                           n6527) );
   NO210  g55( .A(n5580), .B(n5536), .Y(n6528) );
   EN210  g56( .A(n6349), .B(n6348), .Y(n6347) );
   EN210  g57( .A(n6346), .B(n6345), .Y(n6344) );
   EN210  g58( .A(n6343), .B(n6342), .Y(n6341) );
   EN210  g59( .A(n5904), .B(n5907), .Y(n6340) );
   EN210  g60( .A(n5909), .B(n5908), .Y(n5907) );
   BF053  g61( .A1(n5843), .A2(n5842), .B1(n6506), .B2(
                           n6028), .Y(n5689) );
   BF003  g62( .A1(n5687), .A2(n5751), .B1(n5572), .B2(
                           n5689), .Y(n5688) );
   BF053  g63( .A1(n5685), .A2(n5333), .B1(n5573), .B2(
                           n5688), .Y(n5686) );
   BF003  g64( .A1(n5574), .A2(n5686), .B1(n5684), .B2(
                           n5330), .Y(n5575) );
   NO210  g65( .A(n5571), .B(n5328), .Y(n5580) );
   NO210  g66( .A(n6176), .B(n5232), .Y(n5482) );
   NA210  g67( .A(B_6_port), .B(A_12_port), .Y(n5483) );
   NO210  g68( .A(n5652), .B(n5232), .Y(n5484) );
   NA210  g69( .A(B_6_port), .B(A_14_port), .Y(n5910) );
   NO210  g70( .A(n5655), .B(n5232), .Y(n5911) );
   NA210  g71( .A(n5972), .B(n5971), .Y(n6412) );
   NA210  g72( .A(A_2_port), .B(B_2_port), .Y(n6411) );
   NA210  g73( .A(A_3_port), .B(B_1_port), .Y(n5227) );
   NA210  g74( .A(A_5_port), .B(B_0_port), .Y(n5228) );
   NO210  g75( .A(n6478), .B(n5229), .Y(n5455) );
   NA210  g76( .A(B_5_port), .B(A_8_port), .Y(n5979) );
   NA210  g77( .A(A_7_port), .B(B_6_port), .Y(n5980) );
   NA210  g78( .A(A_4_port), .B(B_9_port), .Y(n5981) );
   NO210  g79( .A(n6478), .B(n5982), .Y(n5906) );
   NO210  g80( .A(n6175), .B(n5550), .Y(n5905) );
   NO210  g81( .A(n6478), .B(n6492), .Y(n6252) );
   NO210  g82( .A(n6175), .B(n6070), .Y(n6251) );
   NA210  g83( .A(A_2_port), .B(B_9_port), .Y(n5295) );
   NA210  g84( .A(n5825), .B(n5824), .Y(n5296) );
   NA210  g85( .A(A_3_port), .B(B_8_port), .Y(n6493) );
   NA210  g86( .A(A_4_port), .B(B_11_port), .Y(n6078) );
   NA210  g87( .A(n5837), .B(n5836), .Y(n6137) );
   NA210  g88( .A(A_2_port), .B(B_13_port), .Y(n6136) );
   EN210  g89( .A(n6456), .B(n6014), .Y(n6008) );
   AN210  g90( .A(A_0_port), .B(B_15_port), .Y(n6140) );
   IV110  g91( .A(n5564), .Y(n6300) );
   IV110  g92( .A(n5373), .Y(n5371) );
   IV110  g93( .A(n5563), .Y(n5874) );
   BF053  g94( .A1(n6481), .A2(n6482), .B1(n6441), .B2(
                           n5793), .Y(n6488) );
   IV110  g95( .A(n5562), .Y(n5435) );
   IV110  g96( .A(n5569), .Y(n5955) );
   IV110  g97( .A(n5986), .Y(n5954) );
   IV110  g98( .A(n5994), .Y(n6395) );
   IV110  g99( .A(n5993), .Y(n5873) );
   IV110  g100( .A(n5992), .Y(n5875) );
   EX2B0  g101( .A(n6052), .B(n6094), .Y(n6159) );
   BF053  g102( .A1(n5606), .A2(n6145), .B1(n6081), .B2(
                           n5516), .Y(n5607) );
   EN210  g103( .A(n6149), .B(n6110), .Y(n5756) );
   IV110  g104( .A(n5607), .Y(n5605) );
   EN210  g105( .A(n6581), .B(n6112), .Y(n5332) );
   EN210  g106( .A(n6152), .B(n6539), .Y(n5753) );
   BF003  g107( .A1(n5779), .A2(n6102), .B1(n6516), .B2(
                           n6104), .Y(n5752) );
   EN210  g108( .A(n6155), .B(n6114), .Y(n5750) );
   BF003  g109( .A1(n5778), .A2(n6100), .B1(n6517), .B2(
                           n6101), .Y(n5334) );
   BF003  g110( .A1(n5777), .A2(n6098), .B1(n6518), .B2(
                           n6099), .Y(n5331) );
   IV110  g111( .A(n5434), .Y(n5862) );
   EN210  g112( .A(n5308), .B(n5307), .Y(n5306) );
   BF053  g113( .A1(n6249), .A2(n6248), .B1(n6073), .B2(
                           n5431), .Y(n5863) );
   EN210  g114( .A(n5305), .B(n6263), .Y(n6262) );
   BF053  g115( .A1(n6069), .A2(n5425), .B1(n5865), .B2(
                           n6244), .Y(n5864) );
   IV110  g116( .A(n5864), .Y(n5866) );
   EN2B0  g117( .A(n6424), .B(n6404), .Y(n5734) );
   BF053  g118( .A1(n6072), .A2(n5430), .B1(n6246), .B2(
                           n6245), .Y(n5867) );
   EN210  g119( .A(n5901), .B(n5527), .Y(n5735) );
   IV110  g120( .A(n5867), .Y(n5868) );
   BF053  g121( .A1(n6410), .A2(n6407), .B1(n6411), .B2(
                           n6412), .Y(n6450) );
   BF003  g122( .A1(n6243), .A2(n5966), .B1(n5967), .B2(
                           n6242), .Y(n6451) );
   BF053  g123( .A1(n5343), .A2(n6406), .B1(n6172), .B2(
                           n6451), .Y(n6452) );
   IV110  g124( .A(n6438), .Y(n5349) );
   BF053  g125( .A1(n5225), .A2(n6454), .B1(n6520), .B2(
                           n6519), .Y(n6453) );
   IV110  g126( .A(n6439), .Y(n5348) );
   IV110  g127( .A(n6453), .Y(n6455) );
   IV110  g128( .A(n6441), .Y(n5346) );
   BF053  g129( .A1(n5497), .A2(n5459), .B1(n5230), .B2(
                           n5496), .Y(n5495) );
   IV110  g130( .A(n6443), .Y(n5345) );
   BF051  g131( .A1(n5922), .B1(n5767), .B2(n5942), .Y(
                           n6169) );
   EN2B0  g132( .A(n6172), .B(n6451), .Y(n5343) );
   BF003  g133( .A1(n5886), .A2(n6447), .B1(n5227), .B2(
                           n6015), .Y(n6448) );
   EN2B0  g134( .A(n6413), .B(n6448), .Y(n6519) );
   BF003  g135( .A1(n5885), .A2(n6454), .B1(n5225), .B2(
                           n6452), .Y(n6520) );
   BF003  g136( .A1(n5884), .A2(n6455), .B1(n5228), .B2(
                           n6453), .Y(n5463) );
   IV110  g137( .A(n5664), .Y(n5948) );
   BF003  g138( .A1(n5883), .A2(n5496), .B1(n5230), .B2(
                           n6450), .Y(n5497) );
   IV110  g139( .A(n5662), .Y(n5949) );
   EN210  g140( .A(n5459), .B(n5497), .Y(n5462) );
   IV110  g141( .A(n5928), .Y(n5536) );
   NA210  g142( .A(n6013), .B(n6368), .Y(n5765) );
   IV110  g143( .A(n6516), .Y(n5779) );
   IV110  g144( .A(n6517), .Y(n5778) );
   IV110  g145( .A(n6518), .Y(n5777) );
   EN210  g146( .A(n5301), .B(n6397), .Y(n5903) );
   EN210  g147( .A(n6331), .B(n5935), .Y(n5472) );
   EX210  g148( .A(n5648), .B(n5499), .Y(n5502) );
   EN2B0  g149( .A(n5649), .B(n5501), .Y(n5471) );
   EX210  g150( .A(n6066), .B(n5931), .Y(n6375) );
   NA410  g151( .A(n5926), .B(n6241), .C(n5927), .D(n5928), 
                           .Y(n6361) );
   IV110  g152( .A(n6434), .Y(n5952) );
   BF001  g153( .A1(n5929), .B1(n5583), .B2(n6240), .Y(
                           n5767) );
   IV110  g154( .A(n5481), .Y(n6393) );
   IV110  g155( .A(n5767), .Y(n5769) );
   IV110  g156( .A(n5480), .Y(n5436) );
   BF052  g157( .A1(n6527), .B1(n5945), .B2(n5767), .B3(
                           n5942), .Y(n5341) );
   IV110  g158( .A(n5479), .Y(n5437) );
   NA310  g159( .A(n5928), .B(n6241), .C(n5927), .Y(n6312) );
   IV110  g160( .A(n5477), .Y(n5438) );
   EN210  g161( .A(n6509), .B(n5797), .Y(n6277) );
   BF003  g162( .A1(n5771), .A2(n6531), .B1(n6510), .B2(
                           n6532), .Y(n6276) );
   BF003  g163( .A1(n5770), .A2(n6533), .B1(n6511), .B2(
                           n6535), .Y(n6208) );
   EN210  g164( .A(n6275), .B(n6208), .Y(n6280) );
   BF003  g165( .A1(n5354), .A2(n6536), .B1(n6512), .B2(
                           n6537), .Y(n6279) );
   BF003  g166( .A1(n5911), .A2(n6111), .B1(n5269), .B2(
                           n5624), .Y(n6094) );
   BF053  g167( .A1(n5626), .A2(n5625), .B1(n5660), .B2(
                           n5270), .Y(n5268) );
   IV110  g168( .A(n5268), .Y(n5267) );
   BF053  g169( .A1(n5623), .A2(n5622), .B1(n5919), .B2(
                           n6106), .Y(n5266) );
   IV110  g170( .A(n5266), .Y(n5265) );
   IV110  g171( .A(n5963), .Y(n5961) );
   EX2B0  g172( .A(n6472), .B(n5651), .Y(n5639) );
   BF053  g173( .A1(n6491), .A2(n6287), .B1(n5299), .B2(
                           n5300), .Y(n5960) );
   EN2B0  g174( .A(n5653), .B(n5610), .Y(n5421) );
   IV110  g175( .A(n5960), .Y(n5959) );
   EN210  g176( .A(n5309), .B(n5710), .Y(n5422) );
   BF053  g177( .A1(n6253), .A2(n6250), .B1(n5296), .B2(
                           n5295), .Y(n5958) );
   EX210  g178( .A(n5654), .B(n5713), .Y(n6166) );
   BF053  g179( .A1(n6493), .A2(n5530), .B1(n5956), .B2(
                           n5297), .Y(n5957) );
   BF003  g180( .A1(n6300), .A2(n6116), .B1(n5564), .B2(
                           n6119), .Y(n5848) );
   IV110  g181( .A(n5933), .Y(n5936) );
   EX210  g182( .A(n5554), .B(n5500), .Y(n5930) );
   BF053  g183( .A1(n5403), .A2(n5402), .B1(n5555), .B2(
                           n5504), .Y(n5937) );
   EN210  g184( .A(n5555), .B(n5504), .Y(n5402) );
   BF053  g185( .A1(n5640), .A2(n5936), .B1(n5822), .B2(
                           n5821), .Y(n5938) );
   EN210  g186( .A(n5820), .B(n6375), .Y(n5403) );
   BF053  g187( .A1(n6333), .A2(n6334), .B1(n6335), .B2(
                           n6332), .Y(n5939) );
   EX210  g188( .A(n5556), .B(n5937), .Y(n6377) );
   BF053  g189( .A1(n5641), .A2(n6372), .B1(n6371), .B2(
                           n6338), .Y(n6370) );
   EN210  g190( .A(n5558), .B(n6376), .Y(n5830) );
   NA210  g191( .A(n6330), .B(n5899), .Y(n6334) );
   BF003  g192( .A1(n6392), .A2(n5804), .B1(n5912), .B2(
                           n6109), .Y(n5805) );
   NA210  g193( .A(A_2_port), .B(B_6_port), .Y(n6333) );
   BF003  g194( .A1(n5272), .A2(n6391), .B1(n5273), .B2(
                           n5913), .Y(n6588) );
   NO210  g195( .A(n6478), .B(n5642), .Y(n6337) );
   BF003  g196( .A1(n6390), .A2(n5274), .B1(n5914), .B2(
                           n5690), .Y(n6585) );
   NO210  g197( .A(n6175), .B(n5234), .Y(n6336) );
   BF003  g198( .A1(n6389), .A2(n5691), .B1(n5915), .B2(
                           n5693), .Y(n5808) );
   EN210  g199( .A(n5916), .B(n5808), .Y(n6586) );
   BF003  g200( .A1(n6388), .A2(n5694), .B1(n5917), .B2(
                           n5696), .Y(n6219) );
   IV110  g201( .A(n5535), .Y(n6360) );
   BF003  g202( .A1(n5249), .A2(n5285), .B1(n6076), .B2(
                           n5286), .Y(n6550) );
   IV110  g203( .A(n5926), .Y(n5539) );
   BF003  g204( .A1(n5248), .A2(n6549), .B1(n6084), .B2(
                           n6551), .Y(n5414) );
   IV110  g205( .A(n5940), .Y(n5768) );
   IV110  g206( .A(n6363), .Y(n6294) );
   IV110  g207( .A(n6367), .Y(n5584) );
   IV110  g208( .A(n5587), .Y(n6368) );
   IV110  g209( .A(n6157), .Y(n5759) );
   IV110  g210( .A(n5635), .Y(n5633) );
   NA210  g211( .A(A_0_port), .B(B_2_port), .Y(n5969) );
   NA210  g212( .A(B_1_port), .B(A_1_port), .Y(n5968) );
   NA210  g213( .A(B_0_port), .B(A_3_port), .Y(n6172) );
   NO210  g214( .A(n6478), .B(n6173), .Y(n5972) );
   NO210  g215( .A(n6175), .B(n6174), .Y(n5971) );
   NA210  g216( .A(A_5_port), .B(B_7_port), .Y(n5552) );
   NA210  g217( .A(A_4_port), .B(B_2_port), .Y(n5553) );
   NO210  g218( .A(n5644), .B(n6174), .Y(n5554) );
   NA210  g219( .A(B_2_port), .B(A_6_port), .Y(n5555) );
   NO210  g220( .A(n6174), .B(n5557), .Y(n5556) );
   NA210  g221( .A(A_5_port), .B(B_9_port), .Y(n5235) );
   NA210  g222( .A(B_8_port), .B(A_6_port), .Y(n5236) );
   NA210  g223( .A(A_7_port), .B(B_7_port), .Y(n5237) );
   BF003  g224( .A1(n5347), .A2(n6212), .B1(n6005), .B2(
                           n6214), .Y(n5795) );
   NA210  g225( .A(B_4_port), .B(A_10_port), .Y(n5238) );
   BF003  g226( .A1(n5346), .A2(n5793), .B1(n6441), .B2(
                           n5794), .Y(n6481) );
   NA210  g227( .A(B_0_port), .B(A_6_port), .Y(n5239) );
   EX2B0  g228( .A(n6442), .B(n5792), .Y(n5369) );
   NO210  g229( .A(n6477), .B(n5557), .Y(n5240) );
   BF003  g230( .A1(n5345), .A2(n5374), .B1(n6443), .B2(
                           n5790), .Y(n6065) );
   EN210  g231( .A(n6580), .B(n6579), .Y(n6155) );
   EN210  g232( .A(n5823), .B(n5826), .Y(n5829) );
   EX210  g233( .A(n6583), .B(n6582), .Y(n6581) );
   EN210  g234( .A(n5828), .B(n5827), .Y(n5826) );
   EN210  g235( .A(n5825), .B(n5824), .Y(n5823) );
   EX210  g236( .A(n5822), .B(n5821), .Y(n5820) );
   BF003  g237( .A1(n5244), .A2(n6474), .B1(n5764), .B2(
                           n5733), .Y(n6473) );
   EX210  g238( .A(n5892), .B(n5464), .Y(n5394) );
   BF053  g239( .A1(n5650), .A2(n6473), .B1(n6522), .B2(
                           n6521), .Y(n6472) );
   EX210  g240( .A(n5393), .B(n5392), .Y(n5391) );
   IV110  g241( .A(n5513), .Y(n6556) );
   BF056  g242( .A1(n5255), .A2(n5924), .B1(n5532), .B2(
                           n5580), .Y(n5638) );
   IV110  g243( .A(n6078), .Y(n5254) );
   NA310  g244( .A(n6385), .B(n5258), .C(n6011), .Y(n6215) );
   IV110  g245( .A(n6077), .Y(n5670) );
   IV110  g246( .A(n6083), .Y(n5788) );
   IV110  g247( .A(n5560), .Y(n6302) );
   IV110  g248( .A(n6508), .Y(n6305) );
   IV110  g249( .A(n6507), .Y(n5357) );
   IV110  g250( .A(n6506), .Y(n5364) );
   IV110  g251( .A(n6023), .Y(n6022) );
   BF053  g252( .A1(n5993), .A2(n5278), .B1(n5316), .B2(
                           n5315), .Y(n6021) );
   IV110  g253( .A(n6021), .Y(n6020) );
   BF053  g254( .A1(n5319), .A2(n5318), .B1(n5994), .B2(
                           n5280), .Y(n6019) );
   IV110  g255( .A(n6019), .Y(n6018) );
   BF053  g256( .A1(n6582), .A2(n6583), .B1(n5995), .B2(
                           n5819), .Y(n6017) );
   IV110  g257( .A(n6017), .Y(n6016) );
   BF003  g258( .A1(n6426), .A2(n5818), .B1(n5598), .B2(
                           n5741), .Y(n5599) );
   BF053  g259( .A1(n6427), .A2(n6018), .B1(n5742), .B2(
                           n5743), .Y(n5597) );
   IV110  g260( .A(n5597), .Y(n5596) );
   NA210  g261( .A(A_13_port), .B(B_8_port), .Y(n5912) );
   NA210  g262( .A(B_11_port), .B(A_10_port), .Y(n5913) );
   NA210  g263( .A(A_8_port), .B(B_13_port), .Y(n5914) );
   NA210  g264( .A(A_7_port), .B(B_14_port), .Y(n5915) );
   NA210  g265( .A(A_6_port), .B(B_15_port), .Y(n5916) );
   NA210  g266( .A(B_13_port), .B(A_14_port), .Y(n5487) );
   NA210  g267( .A(A_15_port), .B(B_12_port), .Y(n5488) );
   NA210  g268( .A(n5489), .B(n6480), .Y(n5338) );
   NA210  g269( .A(B_14_port), .B(A_14_port), .Y(n5490) );
   NA210  g270( .A(A_13_port), .B(B_15_port), .Y(n5491) );
   NA210  g271( .A(n5721), .B(n5720), .Y(n5909) );
   NA210  g272( .A(A_2_port), .B(B_11_port), .Y(n5908) );
   NA210  g273( .A(A_3_port), .B(B_10_port), .Y(n5983) );
   NA210  g274( .A(A_5_port), .B(B_8_port), .Y(n5984) );
   NA210  g275( .A(B_7_port), .B(A_6_port), .Y(n5985) );
   NA210  g276( .A(A_5_port), .B(B_12_port), .Y(n5567) );
   NA210  g277( .A(A_7_port), .B(B_10_port), .Y(n5568) );
   NA210  g278( .A(B_7_port), .B(A_10_port), .Y(n5569) );
   NA210  g279( .A(A_11_port), .B(B_7_port), .Y(n5986) );
   NA210  g280( .A(B_8_port), .B(A_10_port), .Y(n5987) );
   IV110  g281( .A(n5758), .Y(n6156) );
   NO210  g282( .A(n6175), .B(n6184), .Y(n6139) );
   IV110  g283( .A(n5632), .Y(n5634) );
   NA210  g284( .A(A_3_port), .B(B_12_port), .Y(n6079) );
   IV110  g285( .A(B_14_port), .Y(n6184) );
   NA210  g286( .A(A_5_port), .B(B_10_port), .Y(n6080) );
   IV110  g287( .A(B_13_port), .Y(n5982) );
   NA210  g288( .A(A_7_port), .B(B_8_port), .Y(n6081) );
   IV110  g289( .A(A_13_port), .Y(n5652) );
   NA210  g290( .A(A_8_port), .B(B_7_port), .Y(n6082) );
   BF053  g291( .A1(n5414), .A2(n5840), .B1(n6084), .B2(
                           n6549), .Y(n6541) );
   BF003  g292( .A1(n5482), .A2(n6541), .B1(n6539), .B2(
                           n6152), .Y(n6540) );
   BF053  g293( .A1(n6114), .A2(n6155), .B1(n5483), .B2(
                           n6540), .Y(n6115) );
   BF003  g294( .A1(n6112), .A2(n6581), .B1(n5484), .B2(
                           n6115), .Y(n6113) );
   BF053  g295( .A1(n6110), .A2(n6149), .B1(n5910), .B2(
                           n6113), .Y(n6111) );
   BF053  g296( .A1(n6108), .A2(n6146), .B1(n6435), .B2(
                           n5599), .Y(n6109) );
   IV110  g297( .A(A_0_port), .Y(n6478) );
   BF053  g298( .A1(n6148), .A2(n6147), .B1(n5481), .B2(
                           n5596), .Y(n6107) );
   IV110  g299( .A(B_2_port), .Y(n6174) );
   IV110  g300( .A(n6107), .Y(n6106) );
   EX2B0  g301( .A(n6425), .B(n6402), .Y(n5611) );
   BF053  g302( .A1(n5826), .A2(n5823), .B1(n5827), .B2(
                           n5828), .Y(n5869) );
   EN2B0  g303( .A(n6177), .B(n5612), .Y(n5737) );
   BF053  g304( .A1(n6071), .A2(n6286), .B1(n6285), .B2(
                           n5829), .Y(n6284) );
   EN210  g305( .A(n5395), .B(n6566), .Y(n5738) );
   BF003  g306( .A1(n6304), .A2(n5711), .B1(n6178), .B2(
                           n6568), .Y(n5710) );
   BF003  g307( .A1(n6303), .A2(n5294), .B1(n5656), .B2(
                           n5712), .Y(n6352) );
   BF003  g308( .A1(n6302), .A2(n6457), .B1(n5560), .B2(
                           n6458), .Y(n5260) );
   EN210  g309( .A(n5844), .B(n5260), .Y(n5998) );
   EN210  g310( .A(n5398), .B(n6290), .Y(n5419) );
   IV110  g311( .A(n5495), .Y(n5498) );
   IV110  g312( .A(n6444), .Y(n6299) );
   BF053  g313( .A1(n5457), .A2(n5458), .B1(n5456), .B2(
                           n6414), .Y(n5499) );
   IV110  g314( .A(n5487), .Y(n6297) );
   BF053  g315( .A1(n5399), .A2(n5400), .B1(n5553), .B2(
                           n5498), .Y(n5500) );
   IV110  g316( .A(n5485), .Y(n6298) );
   BF003  g317( .A1(n5648), .A2(n5499), .B1(n5502), .B2(
                           n5394), .Y(n5501) );
   IV110  g318( .A(n5492), .Y(n6295) );
   IV110  g319( .A(n5490), .Y(n6296) );
   IV110  g320( .A(n6237), .Y(n6382) );
   IV110  g321( .A(n5661), .Y(n5950) );
   BF003  g322( .A1(n5882), .A2(n6449), .B1(n5231), .B2(
                           n6446), .Y(n5461) );
   IV110  g323( .A(n6093), .Y(n6186) );
   BF003  g324( .A1(n5881), .A2(n5718), .B1(n5983), .B2(
                           n6036), .Y(n5719) );
   IV110  g325( .A(n6092), .Y(n6187) );
   IV110  g326( .A(n6091), .Y(n6188) );
   IV110  g327( .A(n6090), .Y(n6189) );
   IV110  g328( .A(n6089), .Y(n6190) );
   IV110  g329( .A(n6087), .Y(n6191) );
   IV110  g340( .A(n6086), .Y(n6192) );
   BF053  g341( .A1(n5383), .A2(n6046), .B1(n5667), .B2(
                           n6223), .Y(n5384) );
   IV110  g342( .A(n5384), .Y(n5382) );
   BF053  g343( .A1(n6048), .A2(n6047), .B1(n5666), .B2(
                           n6221), .Y(n5381) );
   IV110  g344( .A(n5381), .Y(n5380) );
   BF053  g345( .A1(n5378), .A2(n5627), .B1(n5665), .B2(
                           n6218), .Y(n5379) );
   IV110  g346( .A(n5379), .Y(n5377) );
   IV110  g347( .A(n5932), .Y(n6372) );
   BF053  g348( .A1(n5629), .A2(n5628), .B1(n5664), .B2(
                           n6216), .Y(n5376) );
   IV110  g349( .A(n5640), .Y(n5785) );
   IV110  g350( .A(n5376), .Y(n5375) );
   EN2B0  g351( .A(n6067), .B(n6374), .Y(n5474) );
   EN210  g352( .A(n5391), .B(n5432), .Y(n5900) );
   BF003  g353( .A1(n5363), .A2(n5860), .B1(n6068), .B2(
                           n6378), .Y(n5861) );
   BF003  g354( .A1(n5362), .A2(n5862), .B1(n6074), .B2(
                           n5434), .Y(n5902) );
   BF003  g355( .A1(n5361), .A2(n6400), .B1(n6494), .B2(
                           n6401), .Y(n5614) );
   EN210  g356( .A(n5637), .B(n5636), .Y(n6383) );
   EX210  g357( .A(n5534), .B(n5638), .Y(PRODUCT_24_port) );
   EX2B0  g358( .A(n5736), .B(n5639), .Y(PRODUCT_13_port) );
   EN210  g359( .A(n5508), .B(n6056), .Y(PRODUCT_21_port) );
   EX210  g360( .A(n5730), .B(n6057), .Y(PRODUCT_9_port) );
   IV110  g361( .A(n5476), .Y(n5439) );
   IV110  g362( .A(n5475), .Y(n5440) );
   IV110  g363( .A(n6109), .Y(n5804) );
   IV110  g364( .A(n5919), .Y(n6386) );
   IV110  g365( .A(n5918), .Y(n6387) );
   EN210  g366( .A(n5410), .B(n5702), .Y(n5840) );
   EN210  g367( .A(n6344), .B(n6559), .Y(n6349) );
   BF003  g368( .A1(n6201), .A2(n6372), .B1(n5641), .B2(
                           n5932), .Y(n6371) );
   BF003  g369( .A1(n6200), .A2(n6373), .B1(n5647), .B2(
                           n6370), .Y(n5392) );
   EN210  g370( .A(n5390), .B(n5428), .Y(n5393) );
   BF053  g371( .A1(n6224), .A2(n6587), .B1(n5918), .B2(
                           n5697), .Y(n6225) );
   IV110  g372( .A(n6185), .Y(n5454) );
   IV110  g373( .A(n6225), .Y(n6223) );
   IV110  g374( .A(n6079), .Y(n5253) );
   BF053  g375( .A1(n6588), .A2(n5620), .B1(n5913), .B2(
                           n5272), .Y(n6222) );
   IV110  g376( .A(n6500), .Y(n5245) );
   IV110  g377( .A(n6222), .Y(n6221) );
   IV110  g378( .A(n5565), .Y(n5879) );
   BF053  g379( .A1(n5917), .A2(n5694), .B1(n6219), .B2(
                           n6584), .Y(n6220) );
   IV110  g380( .A(n5912), .Y(n6392) );
   BF003  g381( .A1(n5879), .A2(n6234), .B1(n5565), .B2(
                           n6120), .Y(n6235) );
   EN210  g382( .A(n5566), .B(n6235), .Y(n5849) );
   BF003  g383( .A1(n5878), .A2(n6121), .B1(n5567), .B2(
                           n6122), .Y(n6231) );
   BF003  g384( .A1(n5877), .A2(n6230), .B1(n5989), .B2(
                           n6232), .Y(n5812) );
   BF003  g385( .A1(n6233), .A2(n5876), .B1(n5275), .B2(
                           n5990), .Y(n6025) );
   IV110  g386( .A(n5512), .Y(n6465) );
   BF053  g387( .A1(n5235), .A2(n6128), .B1(n6463), .B2(
                           n6256), .Y(n6464) );
   IV110  g388( .A(n6464), .Y(n6462) );
   BF053  g389( .A1(n6181), .A2(n6561), .B1(n6460), .B2(
                           n6262), .Y(n6461) );
   IV110  g390( .A(n6461), .Y(n6459) );
   EN210  g391( .A(n6350), .B(n6578), .Y(n6577) );
   IV110  g392( .A(n6370), .Y(n6373) );
   EN210  g393( .A(n6576), .B(n6575), .Y(n6574) );
   BF003  g394( .A1(n6066), .A2(n5931), .B1(n6375), .B2(
                           n5820), .Y(n6374) );
   EN210  g395( .A(n6573), .B(n6572), .Y(n6571) );
   BF003  g396( .A1(n6377), .A2(n5473), .B1(n5556), .B2(
                           n5937), .Y(n6376) );
   EN210  g397( .A(n6570), .B(n6569), .Y(n6145) );
   BF053  g398( .A1(n5900), .A2(n5474), .B1(n6067), .B2(
                           n6374), .Y(n6378) );
   EN210  g399( .A(n6144), .B(n6143), .Y(n6142) );
   BF053  g400( .A1(n5647), .A2(n6373), .B1(n5393), .B2(
                           n5392), .Y(n6379) );
   BF003  g401( .A1(n5355), .A2(n5526), .B1(n5559), .B2(
                           n5433), .Y(n5527) );
   BF003  g402( .A1(n6309), .A2(n5525), .B1(n5976), .B2(
                           n5528), .Y(n5833) );
   EN210  g403( .A(n5467), .B(n5614), .Y(n5834) );
   BF003  g404( .A1(n6308), .A2(n6470), .B1(n5977), .B2(
                           n6471), .Y(n6566) );
   BF003  g405( .A1(n6307), .A2(n6565), .B1(n6179), .B2(
                           n6567), .Y(n5310) );
   BF003  g406( .A1(n5639), .A2(n5736), .B1(n5651), .B2(
                           n6472), .Y(n5610) );
   BF053  g407( .A1(n5738), .A2(n5737), .B1(n6177), .B2(
                           n5612), .Y(n6568) );
   BF053  g408( .A1(n6566), .A2(n5395), .B1(n5977), .B2(
                           n6470), .Y(n6567) );
   IV110  g409( .A(n6567), .Y(n6565) );
   BF053  g410( .A1(n5397), .A2(n5396), .B1(n6416), .B2(
                           n5613), .Y(n6564) );
   IV110  g411( .A(n5709), .Y(n5707) );
   BF053  g412( .A1(n5705), .A2(n5407), .B1(n6502), .B2(
                           n5603), .Y(n5706) );
   IV110  g413( .A(n5706), .Y(n5704) );
   BF053  g414( .A1(n6504), .A2(n5608), .B1(n5702), .B2(
                           n5410), .Y(n5703) );
   IV110  g415( .A(n5703), .Y(n5701) );
   BF053  g416( .A1(n6154), .A2(n6153), .B1(n5569), .B2(
                           n5701), .Y(n5700) );
   BF003  g417( .A1(n5353), .A2(n6538), .B1(n6513), .B2(
                           n6321), .Y(n6213) );
   IV110  g418( .A(n5700), .Y(n5284) );
   EN210  g419( .A(n6278), .B(n6213), .Y(n6283) );
   BF003  g420( .A1(n5282), .A2(n6267), .B1(n5561), .B2(
                           n6125), .Y(n5283) );
   EN210  g421( .A(n5412), .B(n5411), .Y(n5410) );
   EN210  g422( .A(n5840), .B(n5414), .Y(n5413) );
   EN210  g423( .A(n5843), .B(n5842), .Y(n5841) );
   EN210  g424( .A(n5846), .B(n5845), .Y(n5844) );
   EN210  g425( .A(n5849), .B(n5848), .Y(n5847) );
   EN210  g426( .A(n6266), .B(n6265), .Y(n6264) );
   EX210  g427( .A(n6269), .B(n6268), .Y(n6267) );
   EN210  g428( .A(n5466), .B(n5465), .Y(n5729) );
   EN210  g429( .A(n6272), .B(n6271), .Y(n6270) );
   EN210  g430( .A(n5728), .B(n5727), .Y(n5726) );
   NA210  g431( .A(n5576), .B(n6158), .Y(n5533) );
   BF053  g432( .A1(n5846), .A2(n5845), .B1(n6508), .B2(
                           n6033), .Y(n5683) );
   IV110  g433( .A(n5683), .Y(n5682) );
   BF053  g434( .A1(n5680), .A2(n5841), .B1(n6507), .B2(
                           n6031), .Y(n5681) );
   IV110  g435( .A(n5681), .Y(n5264) );
   BF053  g436( .A1(n5263), .A2(n6163), .B1(n5996), .B2(
                           n5682), .Y(n6000) );
   BF053  g437( .A1(n6164), .A2(n6165), .B1(n5577), .B2(
                           n5264), .Y(n5262) );
   IV110  g438( .A(n5262), .Y(n5261) );
   BF053  g439( .A1(n5260), .A2(n5844), .B1(n5560), .B2(
                           n6457), .Y(n5632) );
   BF053  g440( .A1(n6590), .A2(n6591), .B1(n5578), .B2(
                           n5261), .Y(n5219) );
   NA210  g441( .A(B_2_port), .B(A_8_port), .Y(n5558) );
   NA210  g442( .A(B_2_port), .B(A_9_port), .Y(n5559) );
   NA210  g443( .A(B_2_port), .B(A_10_port), .Y(n5976) );
   NA210  g444( .A(B_2_port), .B(A_11_port), .Y(n5977) );
   NA210  g445( .A(B_4_port), .B(A_9_port), .Y(n5978) );
   NA210  g446( .A(B_4_port), .B(A_12_port), .Y(n6506) );
   NA210  g447( .A(B_3_port), .B(A_13_port), .Y(n6507) );
   NA210  g448( .A(B_2_port), .B(A_14_port), .Y(n6508) );
   NA210  g449( .A(B_1_port), .B(A_15_port), .Y(n5560) );
   NO210  g450( .A(n6423), .B(n5642), .Y(n5561) );
   NA210  g451( .A(n5386), .B(n5385), .Y(n5828) );
   NA210  g452( .A(A_2_port), .B(B_8_port), .Y(n5827) );
   NA210  g453( .A(A_3_port), .B(B_7_port), .Y(n6071) );
   NA210  g454( .A(A_4_port), .B(B_6_port), .Y(n6072) );
   NA210  g455( .A(B_4_port), .B(A_6_port), .Y(n6073) );
   NA210  g456( .A(B_0_port), .B(A_12_port), .Y(n5650) );
   NO210  g457( .A(n6477), .B(n5652), .Y(n5651) );
   NA210  g458( .A(B_0_port), .B(A_14_port), .Y(n5653) );
   EN2B0  g459( .A(n5488), .B(n5370), .Y(n6318) );
   NO210  g460( .A(n6477), .B(n5655), .Y(n5654) );
   NA210  g461( .A(B_0_port), .B(A_8_port), .Y(n5241) );
   BF003  g462( .A1(n6299), .A2(n5371), .B1(n6444), .B2(
                           n5373), .Y(n5365) );
   NO210  g463( .A(n6477), .B(n6423), .Y(n5242) );
   EN210  g464( .A(n6445), .B(n5365), .Y(n6479) );
   NA210  g465( .A(B_0_port), .B(A_10_port), .Y(n5243) );
   EN210  g466( .A(n6064), .B(n5369), .Y(n6482) );
   NO210  g467( .A(n6477), .B(n6176), .Y(n5244) );
   BF003  g468( .A1(n6298), .A2(n6319), .B1(n5485), .B2(
                           n5366), .Y(n6314) );
   EN210  g469( .A(n5486), .B(n6314), .Y(n6485) );
   BF003  g470( .A1(n6297), .A2(n5367), .B1(n5487), .B2(
                           n5368), .Y(n6484) );
   BF053  g471( .A1(n5834), .A2(n5833), .B1(n5976), .B2(
                           n5525), .Y(n6471) );
   EN210  g472( .A(n6339), .B(n5387), .Y(n5390) );
   IV110  g473( .A(n6471), .Y(n6470) );
   EN210  g474( .A(n5389), .B(n5388), .Y(n5387) );
   BF053  g475( .A1(n5468), .A2(n5469), .B1(n6495), .B2(
                           n6396), .Y(n6469) );
   IV110  g476( .A(n6469), .Y(n6468) );
   BF003  g477( .A1(n5443), .A2(n6024), .B1(n6430), .B2(
                           n5810), .Y(n5590) );
   BF053  g478( .A1(n6045), .A2(n5729), .B1(n6496), .B2(
                           n5964), .Y(n6467) );
   EN210  g479( .A(n6431), .B(n5590), .Y(n5322) );
   IV110  g480( .A(n6467), .Y(n6044) );
   BF003  g481( .A1(n5449), .A2(n5529), .B1(n6498), .B2(
                           n5957), .Y(n5727) );
   BF003  g482( .A1(n5448), .A2(n6037), .B1(n5984), .B2(
                           n6038), .Y(n6131) );
   BF003  g483( .A1(n5447), .A2(n6130), .B1(n5236), .B2(
                           n6132), .Y(n6260) );
   BF003  g484( .A1(n5446), .A2(n6286), .B1(n6071), .B2(
                           n5426), .Y(n6285) );
   EN210  g485( .A(n5297), .B(n5956), .Y(n5300) );
   BF003  g486( .A1(n5445), .A2(n6287), .B1(n6491), .B2(
                           n6284), .Y(n5299) );
   BF003  g487( .A1(n5679), .A2(n5959), .B1(n5552), .B2(
                           n5960), .Y(n6040) );
   BF003  g488( .A1(n5678), .A2(n6039), .B1(n5985), .B2(
                           n6041), .Y(n6345) );
   EN210  g489( .A(n6341), .B(n6131), .Y(n6346) );
   BF003  g490( .A1(n5677), .A2(n6133), .B1(n5237), .B2(
                           n6134), .Y(n5519) );
   IV110  g491( .A(n6535), .Y(n6533) );
   BF053  g492( .A1(n5851), .A2(n5850), .B1(n6089), .B2(
                           n5375), .Y(n6532) );
   IV110  g493( .A(n6532), .Y(n6531) );
   BF053  g494( .A1(n6088), .A2(n6529), .B1(n6087), .B2(
                           n6327), .Y(n6530) );
   IV110  g495( .A(n6530), .Y(n6105) );
   NO210  g496( .A(n5945), .B(n5944), .Y(n5943) );
   NA210  g497( .A(n6515), .B(n5325), .Y(n5928) );
   NO210  g498( .A(n5942), .B(n5941), .Y(n5940) );
   BF053  g499( .A1(n6103), .A2(n5413), .B1(n6505), .B2(
                           n6026), .Y(n6104) );
   NA210  g500( .A(n5510), .B(n5509), .Y(n5508) );
   NA210  g501( .A(A_15_port), .B(B_13_port), .Y(n5492) );
   NA210  g502( .A(n6488), .B(n6487), .Y(n5545) );
   OR210  g503( .A(n6486), .B(n5338), .Y(n5493) );
   NA210  g504( .A(n5548), .B(n5547), .Y(n5336) );
   NO210  g505( .A(n5335), .B(n5336), .Y(n5494) );
   EN210  g506( .A(n5409), .B(n5408), .Y(n5407) );
   EN210  g507( .A(n5406), .B(n5405), .Y(n6359) );
   EN210  g508( .A(n6358), .B(n6354), .Y(n6357) );
   EN210  g509( .A(n6356), .B(n6355), .Y(n6354) );
   EX210  g510( .A(n6353), .B(n6352), .Y(n6351) );
   NA210  g511( .A(A_8_port), .B(B_10_port), .Y(n5988) );
   NA210  g512( .A(A_6_port), .B(B_12_port), .Y(n5989) );
   NA210  g513( .A(A_4_port), .B(B_14_port), .Y(n5990) );
   NA210  g514( .A(A_3_port), .B(B_15_port), .Y(n5991) );
   NA210  g515( .A(A_5_port), .B(B_13_port), .Y(n5992) );
   NO210  g516( .A(n5575), .B(n5754), .Y(n6162) );
   NA210  g517( .A(n5757), .B(n6162), .Y(n5576) );
   NO210  g518( .A(n6158), .B(n5576), .Y(n6241) );
   NA210  g519( .A(B_3_port), .B(A_14_port), .Y(n5577) );
   NA210  g520( .A(B_3_port), .B(A_15_port), .Y(n5578) );
   IV110  g521( .A(A_11_port), .Y(n6176) );
   NA210  g522( .A(B_5_port), .B(A_10_port), .Y(n6083) );
   IV110  g523( .A(B_5_port), .Y(n5229) );
   IV110  g524( .A(B_9_port), .Y(n5646) );
   IV110  g525( .A(B_10_port), .Y(n6070) );
   NA210  g526( .A(B_10_port), .B(A_12_port), .Y(n5667) );
   NA210  g527( .A(A_13_port), .B(B_9_port), .Y(n5668) );
   NA210  g528( .A(A_15_port), .B(B_7_port), .Y(n5669) );
   IV110  g529( .A(n5958), .Y(n5618) );
   NA210  g530( .A(B_9_port), .B(A_14_port), .Y(n6086) );
   IV110  g531( .A(A_15_port), .Y(n5655) );
   BF053  g532( .A1(n5698), .A2(n5747), .B1(n5475), .B2(
                           n6542), .Y(n5699) );
   IV110  g533( .A(B_11_port), .Y(n6492) );
   IV110  g534( .A(n5699), .Y(n5697) );
   IV110  g535( .A(B_3_port), .Y(n6173) );
   IV110  g536( .A(B_12_port), .Y(n5550) );
   IV110  g537( .A(n5225), .Y(n5885) );
   IV110  g538( .A(n5227), .Y(n5886) );
   IV110  g539( .A(n5230), .Y(n5883) );
   IV110  g540( .A(n5233), .Y(n5786) );
   IV110  g541( .A(n5716), .Y(n5714) );
   BF053  g542( .A1(n5422), .A2(n5421), .B1(n5653), .B2(
                           n5610), .Y(n5713) );
   BF053  g543( .A1(n5710), .A2(n5309), .B1(n6178), .B2(
                           n5711), .Y(n5712) );
   IV110  g544( .A(n5712), .Y(n5294) );
   BF053  g545( .A1(n5310), .A2(n5311), .B1(n6179), .B2(
                           n6565), .Y(n5293) );
   IV110  g546( .A(n5293), .Y(n5292) );
   BF003  g547( .A1(n5953), .A2(n5819), .B1(n5995), .B2(
                           n6226), .Y(n6582) );
   BF053  g548( .A1(n5290), .A2(n5306), .B1(n6180), .B2(
                           n6563), .Y(n5291) );
   EN210  g549( .A(n6146), .B(n6108), .Y(n6151) );
   IV110  g550( .A(n5291), .Y(n5289) );
   BF053  g551( .A1(n5552), .A2(n5959), .B1(n6040), .B2(
                           n5726), .Y(n6041) );
   IV110  g552( .A(n6041), .Y(n6039) );
   BF053  g553( .A1(n6498), .A2(n5529), .B1(n5727), .B2(
                           n5728), .Y(n6038) );
   IV110  g554( .A(n6038), .Y(n6037) );
   BF053  g555( .A1(n5723), .A2(n5724), .B1(n5722), .B2(
                           n5304), .Y(n6036) );
   BF053  g556( .A1(n5617), .A2(n5725), .B1(n5551), .B2(
                           n5618), .Y(n5619) );
   IV110  g557( .A(n5619), .Y(n5616) );
   BF053  g558( .A1(n6494), .A2(n6400), .B1(n5614), .B2(
                           n5467), .Y(n5615) );
   IV110  g559( .A(n5615), .Y(n5613) );
   BF003  g560( .A1(n6425), .A2(n6402), .B1(n5611), .B2(
                           n5832), .Y(n5612) );
   EN2B0  g561( .A(n6073), .B(n5431), .Y(n6248) );
   EN210  g562( .A(n6244), .B(n5865), .Y(n6249) );
   BF003  g563( .A1(n5784), .A2(n6398), .B1(n6075), .B2(
                           n5863), .Y(n6397) );
   BF003  g564( .A1(n5783), .A2(n6396), .B1(n6495), .B2(
                           n6399), .Y(n5468) );
   BF003  g565( .A1(n5782), .A2(n6468), .B1(n5978), .B2(
                           n6469), .Y(n5715) );
   BF003  g566( .A1(n5781), .A2(n5714), .B1(n5238), .B2(
                           n5716), .Y(n5307) );
   EN210  g567( .A(n6262), .B(n6460), .Y(n5308) );
   BF003  g568( .A1(n5780), .A2(n5287), .B1(n5659), .B2(
                           n5288), .Y(n6029) );
   BF003  g569( .A1(n5364), .A2(n6028), .B1(n6506), .B2(
                           n6030), .Y(n5842) );
   EN210  g570( .A(n6574), .B(n6029), .Y(n6350) );
   IV110  g571( .A(n5939), .Y(n5429) );
   BF053  g572( .A1(n5663), .A2(n6328), .B1(n5662), .B2(
                           n5807), .Y(n6329) );
   IV110  g573( .A(n5647), .Y(n6200) );
   IV110  g574( .A(n6329), .Y(n6327) );
   IV110  g575( .A(n6378), .Y(n5860) );
   IV110  g576( .A(n6069), .Y(n6199) );
   IV110  g577( .A(n5426), .Y(n6286) );
   IV110  g578( .A(n6072), .Y(n5675) );
   IV110  g579( .A(n5433), .Y(n5526) );
   IV110  g580( .A(n6074), .Y(n5362) );
   EN210  g581( .A(n6060), .B(n6059), .Y(n6058) );
   EN210  g582( .A(n6063), .B(n6062), .Y(n6061) );
   EX210  g583( .A(n6479), .B(n6065), .Y(n6064) );
   EX210  g584( .A(n6482), .B(n6481), .Y(n6480) );
   EN210  g585( .A(n6485), .B(n6484), .Y(n6483) );
   NA210  g586( .A(B_3_port), .B(A_6_port), .Y(n6067) );
   NA210  g587( .A(B_3_port), .B(A_7_port), .Y(n6068) );
   NA210  g588( .A(A_5_port), .B(B_5_port), .Y(n6069) );
   NO210  g589( .A(n6478), .B(n6070), .Y(n5825) );
   NO210  g590( .A(n6175), .B(n5646), .Y(n5824) );
   BF003  g591( .A1(n6199), .A2(n5425), .B1(n6069), .B2(
                           n6379), .Y(n5865) );
   EN210  g592( .A(n5298), .B(n5962), .Y(n5303) );
   BF003  g593( .A1(n6198), .A2(n5866), .B1(n6489), .B2(
                           n5864), .Y(n5302) );
   BF003  g594( .A1(n6197), .A2(n5964), .B1(n6496), .B2(
                           n5965), .Y(n6045) );
   BF003  g595( .A1(n6196), .A2(n6044), .B1(n5979), .B2(
                           n6467), .Y(n6348) );
   EN210  g596( .A(n6586), .B(n6585), .Y(n6584) );
   EN210  g597( .A(n5620), .B(n6588), .Y(n6587) );
   EN210  g598( .A(n5623), .B(n5622), .Y(n5621) );
   EX210  g599( .A(n5626), .B(n5625), .Y(n5624) );
   EN210  g600( .A(n5629), .B(n5628), .Y(n5627) );
   IV110  g601( .A(n6241), .Y(n5532) );
   IV110  g602( .A(n6002), .Y(n5506) );
   IV110  g603( .A(n6004), .Y(n6012) );
   IV110  g604( .A(n5922), .Y(n5941) );
   IV110  g605( .A(n5924), .Y(n6526) );
   BF056  g606( .A1(n6215), .A2(n6002), .B1(n6012), .B2(
                           n5507), .Y(n6056) );
   BF053  g607( .A1(n6213), .A2(n6278), .B1(n6513), .B2(
                           n6538), .Y(n6214) );
   IV110  g608( .A(n6214), .Y(n6212) );
   BF053  g609( .A1(n6280), .A2(n6279), .B1(n6512), .B2(
                           n6536), .Y(n6211) );
   IV110  g610( .A(n6211), .Y(n6210) );
   BF003  g611( .A1(n5654), .A2(n5713), .B1(n6166), .B2(
                           n6351), .Y(n5999) );
   BF003  g612( .A1(n6193), .A2(n5267), .B1(n5669), .B2(
                           n5268), .Y(n6053) );
   BF053  g613( .A1(n6352), .A2(n6353), .B1(n5656), .B2(
                           n5294), .Y(n6458) );
   BF003  g614( .A1(n6192), .A2(n6325), .B1(n6086), .B2(
                           n6326), .Y(n5856) );
   IV110  g615( .A(n6458), .Y(n6457) );
   BF003  g616( .A1(n6191), .A2(n6327), .B1(n6087), .B2(
                           n6329), .Y(n6529) );
   BF053  g617( .A1(n5657), .A2(n5292), .B1(n6034), .B2(
                           n6577), .Y(n6035) );
   EN210  g618( .A(n6088), .B(n6529), .Y(n5851) );
   IV110  g619( .A(n6035), .Y(n6033) );
   BF003  g620( .A1(n6190), .A2(n5375), .B1(n6089), .B2(
                           n5376), .Y(n5850) );
   IV110  g621( .A(n6379), .Y(n5425) );
   BF003  g622( .A1(n6306), .A2(n5292), .B1(n5657), .B2(
                           n5293), .Y(n6034) );
   BF053  g623( .A1(n5387), .A2(n6339), .B1(n5388), .B2(
                           n5389), .Y(n5426) );
   BF003  g624( .A1(n6305), .A2(n6033), .B1(n6508), .B2(
                           n6035), .Y(n5845) );
   BF053  g625( .A1(n5645), .A2(n5429), .B1(n5428), .B2(
                           n5390), .Y(n5427) );
   EN210  g626( .A(n6577), .B(n6034), .Y(n6353) );
   IV110  g627( .A(n5427), .Y(n5430) );
   EN210  g628( .A(n5473), .B(n6377), .Y(n5732) );
   BF003  g629( .A1(n5643), .A2(n5938), .B1(n5432), .B2(
                           n5391), .Y(n5431) );
   EX2B0  g630( .A(n6417), .B(n6288), .Y(n6290) );
   BF003  g631( .A1(n5352), .A2(n6322), .B1(n6514), .B2(
                           n6323), .Y(n6282) );
   BF053  g632( .A1(n5562), .A2(n5704), .B1(n6268), .B2(
                           n6269), .Y(n5281) );
   EN210  g633( .A(n6281), .B(n5920), .Y(n5326) );
   IV110  g634( .A(n5281), .Y(n5280) );
   BF003  g635( .A1(n5351), .A2(n6210), .B1(n6436), .B2(
                           n6211), .Y(n6062) );
   BF003  g636( .A1(n5350), .A2(n6207), .B1(n6437), .B2(
                           n6209), .Y(n5791) );
   BF003  g637( .A1(n5349), .A2(n5799), .B1(n6438), .B2(
                           n6206), .Y(n6059) );
   BF003  g638( .A1(n5348), .A2(n5796), .B1(n6439), .B2(
                           n5798), .Y(n5372) );
   EN210  g639( .A(n6440), .B(n5372), .Y(n6060) );
   EN210  g640( .A(n6058), .B(n5791), .Y(n6063) );
   EN210  g641( .A(n5316), .B(n5315), .Y(n6273) );
   EN210  g642( .A(n5304), .B(n5722), .Y(n5725) );
   EN210  g643( .A(n5319), .B(n5318), .Y(n5317) );
   EN210  g644( .A(n5724), .B(n5723), .Y(n5722) );
   EN210  g645( .A(n5721), .B(n5720), .Y(n5304) );
   EN210  g646( .A(n5303), .B(n5302), .Y(n5301) );
   IV110  g647( .A(n5957), .Y(n5529) );
   EN210  g648( .A(n5300), .B(n5299), .Y(n5298) );
   BF053  g649( .A1(n5559), .A2(n5526), .B1(n5527), .B2(
                           n5901), .Y(n5528) );
   EN210  g650( .A(n6250), .B(n6253), .Y(n5297) );
   BF003  g651( .A1(n5880), .A2(n5717), .B1(n6183), .B2(
                           n6126), .Y(n6257) );
   BF003  g652( .A1(n5454), .A2(n6466), .B1(n6185), .B2(
                           n6127), .Y(n5511) );
   EN210  g653( .A(n6255), .B(n5511), .Y(n6258) );
   BF003  g654( .A1(n5453), .A2(n5618), .B1(n5551), .B2(
                           n5958), .Y(n5617) );
   EN210  g655( .A(n6340), .B(n5719), .Y(n6343) );
   BF003  g656( .A1(n5452), .A2(n5616), .B1(n5981), .B2(
                           n5619), .Y(n6342) );
   BF003  g657( .A1(n5451), .A2(n6128), .B1(n5235), .B2(
                           n6129), .Y(n6463) );
   EN210  g658( .A(n6256), .B(n6463), .Y(n6261) );
   BF003  g659( .A1(n5450), .A2(n5530), .B1(n6493), .B2(
                           n5869), .Y(n5956) );
   EN210  g660( .A(n5725), .B(n5617), .Y(n5728) );
   NA210  g661( .A(A_8_port), .B(B_9_port), .Y(n5562) );
   NA210  g662( .A(A_6_port), .B(B_11_port), .Y(n5563) );
   NA210  g663( .A(A_4_port), .B(B_13_port), .Y(n5564) );
   NA210  g664( .A(A_3_port), .B(B_14_port), .Y(n5565) );
   NA210  g665( .A(A_2_port), .B(B_15_port), .Y(n5566) );
   NA210  g666( .A(n5858), .B(n5329), .Y(n6515) );
   NA210  g667( .A(B_5_port), .B(A_12_port), .Y(n6516) );
   NA210  g668( .A(B_5_port), .B(A_13_port), .Y(n6517) );
   IV110  g669( .A(n5235), .Y(n5451) );
   NA210  g670( .A(B_5_port), .B(A_14_port), .Y(n6518) );
   EX2B0  g671( .A(n6483), .B(n6318), .Y(n6487) );
   NA210  g672( .A(B_1_port), .B(A_14_port), .Y(n5656) );
   EN210  g673( .A(n6480), .B(n5489), .Y(n5335) );
   NA210  g674( .A(B_2_port), .B(A_13_port), .Y(n5657) );
   EX2B0  g675( .A(n6061), .B(n5795), .Y(n5547) );
   NA210  g676( .A(B_3_port), .B(A_12_port), .Y(n5658) );
   BF003  g677( .A1(n6296), .A2(n6313), .B1(n5490), .B2(
                           n6315), .Y(n6310) );
   NA210  g678( .A(B_4_port), .B(A_11_port), .Y(n5659) );
   EN210  g679( .A(n5491), .B(n6310), .Y(n5542) );
   NA210  g680( .A(A_9_port), .B(B_6_port), .Y(n6076) );
   BF003  g681( .A1(n5442), .A2(n5811), .B1(n6432), .B2(
                           n5813), .Y(n6546) );
   BF053  g682( .A1(n6497), .A2(n5961), .B1(n5465), .B2(
                           n5466), .Y(n6043) );
   EN210  g683( .A(n5320), .B(n6546), .Y(n5740) );
   IV110  g684( .A(n6043), .Y(n6042) );
   BF003  g685( .A1(n5441), .A2(n5814), .B1(n6433), .B2(
                           n5816), .Y(n6543) );
   BF003  g686( .A1(n5440), .A2(n6542), .B1(n5475), .B2(
                           n6544), .Y(n5698) );
   BF003  g687( .A1(n5439), .A2(n6545), .B1(n5476), .B2(
                           n6547), .Y(n5695) );
   BF003  g688( .A1(n5438), .A2(n6548), .B1(n5477), .B2(
                           n5591), .Y(n5692) );
   EN210  g689( .A(n5478), .B(n5692), .Y(n5746) );
   BF003  g690( .A1(n5437), .A2(n5592), .B1(n5479), .B2(
                           n5593), .Y(n5745) );
   AN210  g691( .A(n6365), .B(n5540), .Y(n5763) );
   NO210  g692( .A(n5544), .B(n5545), .Y(n6366) );
   NA410  g693( .A(n6369), .B(n6368), .C(n5415), .D(n6237), 
                           .Y(n6367) );
   NO210  g694( .A(n5543), .B(n5493), .Y(n6381) );
   NA210  g695( .A(n5337), .B(n5494), .Y(n5416) );
   EX2B0  g696( .A(n5998), .B(n5999), .Y(PRODUCT_16_port) );
   EX2B0  g697( .A(n5967), .B(n6242), .Y(PRODUCT_2_port) );
   EX210  g698( .A(n5418), .B(n5417), .Y(PRODUCT_10_port) );
   EX2B0  g699( .A(n5420), .B(n5419), .Y(PRODUCT_6_port) );
   EX2B0  g700( .A(n5631), .B(n5997), .Y(PRODUCT_17_port) );
   IV110  g701( .A(n6104), .Y(n6102) );
   NO210  g702( .A(n5507), .B(n5506), .Y(n5505) );
   BF053  g703( .A1(n5752), .A2(n5753), .B1(n6516), .B2(
                           n6102), .Y(n6101) );
   NA210  g704( .A(B_15_port), .B(A_15_port), .Y(n6456) );
   IV110  g705( .A(n6101), .Y(n6100) );
   NA210  g706( .A(B_2_port), .B(A_12_port), .Y(n6179) );
   NA210  g707( .A(B_3_port), .B(A_11_port), .Y(n6180) );
   NA210  g708( .A(B_5_port), .B(A_9_port), .Y(n6181) );
   NA210  g709( .A(A_8_port), .B(B_6_port), .Y(n6182) );
   NA210  g710( .A(A_4_port), .B(B_10_port), .Y(n6183) );
   NA210  g711( .A(n5219), .B(n5220), .Y(n5222) );
   NO210  g712( .A(n5223), .B(n5222), .Y(n5579) );
   NA210  g713( .A(B_2_port), .B(A_15_port), .Y(n5996) );
   NO210  g714( .A(n5999), .B(n5998), .Y(n5997) );
   NO210  g715( .A(n5634), .B(n5635), .Y(n5637) );
   NA210  g716( .A(n5762), .B(n6366), .Y(n6013) );
   NA210  g717( .A(n5760), .B(n5761), .Y(n6014) );
   NA210  g718( .A(n5344), .B(n5763), .Y(n6007) );
   IV110  g719( .A(n5570), .Y(n5776) );
   NO210  g720( .A(n5339), .B(n5923), .Y(n5538) );
   IV110  g721( .A(n6498), .Y(n5449) );
   NA210  g722( .A(A_9_port), .B(B_14_port), .Y(n6087) );
   IV110  g723( .A(n5976), .Y(n6309) );
   NA210  g724( .A(A_8_port), .B(B_15_port), .Y(n6088) );
   IV110  g725( .A(n5239), .Y(n6301) );
   NA210  g726( .A(A_10_port), .B(B_13_port), .Y(n6089) );
   IV110  g727( .A(n5977), .Y(n6308) );
   NA210  g728( .A(A_11_port), .B(B_12_port), .Y(n6090) );
   IV110  g729( .A(n5978), .Y(n5782) );
   NA210  g730( .A(B_11_port), .B(A_12_port), .Y(n6091) );
   BF003  g731( .A1(n5952), .A2(n6016), .B1(n6434), .B2(
                           n6017), .Y(n6150) );
   BF053  g732( .A1(n5308), .A2(n5307), .B1(n5238), .B2(
                           n5714), .Y(n5288) );
   BF003  g733( .A1(n5951), .A2(n5270), .B1(n5660), .B2(
                           n5271), .Y(n5625) );
   IV110  g734( .A(n5288), .Y(n5287) );
   EX2B0  g735( .A(n5482), .B(n6541), .Y(n6539) );
   EN2B0  g736( .A(n5483), .B(n6540), .Y(n6114) );
   EX2B0  g737( .A(n5484), .B(n6115), .Y(n6112) );
   EN2B0  g738( .A(n5910), .B(n6113), .Y(n6110) );
   EX2B0  g739( .A(n5911), .B(n6111), .Y(n5269) );
   BF003  g740( .A1(n5950), .A2(n5803), .B1(n5661), .B2(
                           n5806), .Y(n5801) );
   EN210  g741( .A(n5531), .B(n6240), .Y(PRODUCT_22_port) );
   EX210  g742( .A(n5761), .B(n5760), .Y(n5344) );
   EX2B0  g743( .A(n5344), .B(n5763), .Y(n5762) );
   EX2B0  g744( .A(n5733), .B(n5764), .Y(PRODUCT_11_port) );
   EX2B0  g745( .A(n6236), .B(n5765), .Y(PRODUCT_29_port) );
   EX210  g746( .A(n5312), .B(n5766), .Y(PRODUCT_7_port) );
   BF003  g747( .A1(n5768), .A2(n5767), .B1(n5940), .B2(
                           n5769), .Y(PRODUCT_26_port) );
   EX2B0  g748( .A(n6351), .B(n6166), .Y(PRODUCT_15_port) );
   EX2B0  g749( .A(n6239), .B(n6167), .Y(PRODUCT_23_port) );
   EN210  g750( .A(n5505), .B(n6168), .Y(PRODUCT_20_port) );
   EN210  g751( .A(n5756), .B(n5755), .Y(n5754) );
   BF003  g752( .A1(n5759), .A2(n5758), .B1(n6157), .B2(
                           n6156), .Y(n5757) );
   EN210  g753( .A(n6160), .B(n6159), .Y(n6158) );
   EX210  g754( .A(n6162), .B(n5757), .Y(n6161) );
   EN210  g755( .A(n6165), .B(n6164), .Y(n6163) );
   EX210  g756( .A(n6591), .B(n6590), .Y(n6589) );
   EN210  g757( .A(n5220), .B(n5219), .Y(n6592) );
   EX2B0  g758( .A(n5969), .B(n5968), .Y(n5967) );
   EX210  g759( .A(n5223), .B(n5222), .Y(n5221) );
   EX2B0  g760( .A(n5966), .B(n6243), .Y(n6242) );
   BF003  g761( .A1(n6442), .A2(n5792), .B1(n5369), .B2(
                           n6064), .Y(n5370) );
   BF053  g762( .A1(n6065), .A2(n6479), .B1(n6443), .B2(
                           n5374), .Y(n5368) );
   IV110  g763( .A(n5368), .Y(n5367) );
   BF053  g764( .A1(n6445), .A2(n5365), .B1(n6444), .B2(
                           n5371), .Y(n5366) );
   IV110  g765( .A(n5366), .Y(n6319) );
   BF053  g766( .A1(n6318), .A2(n6483), .B1(n5488), .B2(
                           n5370), .Y(n6365) );
   IV110  g767( .A(n5990), .Y(n5876) );
   BF053  g768( .A1(n6485), .A2(n6484), .B1(n5487), .B2(
                           n5367), .Y(n6317) );
   IV110  g769( .A(n5989), .Y(n5877) );
   IV110  g770( .A(n6317), .Y(n6316) );
   EX2B0  g771( .A(n5572), .B(n5689), .Y(n5687) );
   IV110  g772( .A(n6554), .Y(n6552) );
   EN2B0  g773( .A(n5573), .B(n5688), .Y(n5685) );
   BF053  g774( .A1(n6076), .A2(n5285), .B1(n6550), .B2(
                           n6571), .Y(n6551) );
   EX2B0  g775( .A(n5574), .B(n5686), .Y(n5684) );
   EN210  g776( .A(n5575), .B(n5754), .Y(n5223) );
   EN210  g777( .A(n5333), .B(n5685), .Y(n6591) );
   EN210  g778( .A(n5751), .B(n5687), .Y(n6165) );
   BF003  g779( .A1(n5775), .A2(n5264), .B1(n5577), .B2(
                           n5681), .Y(n6164) );
   BF003  g780( .A1(n5774), .A2(n5261), .B1(n5578), .B2(
                           n5262), .Y(n6590) );
   EN210  g781( .A(n6048), .B(n6047), .Y(n6046) );
   EN210  g782( .A(n6051), .B(n6050), .Y(n6049) );
   EN210  g783( .A(n5386), .B(n5385), .Y(n6339) );
   EN210  g784( .A(n6054), .B(n6053), .Y(n6052) );
   EN210  g785( .A(n6335), .B(n6332), .Y(n6338) );
   EN210  g786( .A(n5851), .B(n5850), .Y(n6055) );
   EN210  g787( .A(n6337), .B(n6336), .Y(n6335) );
   EN210  g788( .A(n5854), .B(n5853), .Y(n5852) );
   EN210  g789( .A(n6334), .B(n6333), .Y(n6332) );
   EN210  g790( .A(n5898), .B(n5895), .Y(n6331) );
   BF053  g791( .A1(n6208), .A2(n6275), .B1(n6511), .B2(
                           n6533), .Y(n6209) );
   IV110  g792( .A(n6505), .Y(n5787) );
   IV110  g793( .A(n6209), .Y(n6207) );
   IV110  g794( .A(n6504), .Y(n6202) );
   BF053  g795( .A1(n6277), .A2(n6276), .B1(n6510), .B2(
                           n6531), .Y(n6206) );
   IV110  g796( .A(n6503), .Y(n6203) );
   IV110  g797( .A(n6206), .Y(n5799) );
   IV110  g798( .A(n6502), .Y(n6204) );
   BF053  g799( .A1(n6509), .A2(n5797), .B1(n6095), .B2(
                           n6105), .Y(n5798) );
   IV110  g800( .A(n6501), .Y(n6205) );
   BF003  g801( .A1(n6189), .A2(n5377), .B1(n6090), .B2(
                           n5379), .Y(n6534) );
   EN210  g802( .A(n6055), .B(n6534), .Y(n5854) );
   BF003  g803( .A1(n6188), .A2(n5380), .B1(n6091), .B2(
                           n5381), .Y(n5853) );
   BF003  g804( .A1(n6187), .A2(n5382), .B1(n6092), .B2(
                           n5384), .Y(n6320) );
   EN210  g805( .A(n5852), .B(n6320), .Y(n5857) );
   BF053  g806( .A1(n5324), .A2(n5740), .B1(n6428), .B2(
                           n6020), .Y(n5595) );
   IV110  g807( .A(n5595), .Y(n5594) );
   BF053  g808( .A1(n6429), .A2(n6022), .B1(n5321), .B2(
                           n5322), .Y(n5593) );
   IV110  g809( .A(n5593), .Y(n5592) );
   BF053  g810( .A1(n6431), .A2(n5590), .B1(n6430), .B2(
                           n6024), .Y(n5591) );
   EN2B0  g811( .A(n6419), .B(n6289), .Y(n5313) );
   EN210  g812( .A(n5470), .B(n5930), .Y(n5314) );
   EX2B0  g813( .A(n6420), .B(n6291), .Y(n6293) );
   EN2B0  g814( .A(n6421), .B(n6292), .Y(n5731) );
   EX2B0  g815( .A(n6422), .B(n6405), .Y(n6403) );
   BF053  g816( .A1(n5985), .A2(n6039), .B1(n6346), .B2(
                           n6345), .Y(n6134) );
   IV110  g817( .A(n6134), .Y(n6133) );
   BF053  g818( .A1(n5984), .A2(n6037), .B1(n6131), .B2(
                           n6341), .Y(n6132) );
   IV110  g819( .A(n6132), .Y(n6130) );
   BF053  g820( .A1(n5981), .A2(n5616), .B1(n6342), .B2(
                           n6343), .Y(n6129) );
   IV110  g821( .A(n5507), .Y(n5258) );
   IV110  g822( .A(n6446), .Y(n6449) );
   IV110  g823( .A(n6005), .Y(n5347) );
   IV110  g824( .A(n6436), .Y(n5351) );
   IV110  g825( .A(n6437), .Y(n5350) );
   BF003  g826( .A1(n5360), .A2(n5613), .B1(n6416), .B2(
                           n5615), .Y(n5396) );
   EN210  g827( .A(n6347), .B(n5715), .Y(n5397) );
   BF003  g828( .A1(n5359), .A2(n6563), .B1(n6180), .B2(
                           n6564), .Y(n5290) );
   BF003  g829( .A1(n5358), .A2(n5289), .B1(n5658), .B2(
                           n5291), .Y(n6578) );
   BF003  g830( .A1(n5357), .A2(n6031), .B1(n6507), .B2(
                           n6032), .Y(n5680) );
   IV110  g831( .A(n6220), .Y(n6218) );
   BF053  g832( .A1(n5914), .A2(n5274), .B1(n6585), .B2(
                           n6586), .Y(n6217) );
   IV110  g833( .A(n6217), .Y(n6216) );
   BF053  g834( .A1(n5915), .A2(n5691), .B1(n5916), .B2(
                           n5808), .Y(n5809) );
   IV110  g835( .A(n5809), .Y(n5807) );
   BF053  g836( .A1(n5912), .A2(n5804), .B1(n5805), .B2(
                           n5621), .Y(n5806) );
   IV110  g837( .A(n6381), .Y(n5888) );
   IV110  g838( .A(n5806), .Y(n5803) );
   IV110  g839( .A(n5416), .Y(n5944) );
   BF053  g840( .A1(n6054), .A2(n6053), .B1(n5669), .B2(
                           n5267), .Y(n5859) );
   IV110  g841( .A(n5528), .Y(n5525) );
   EN210  g842( .A(n5296), .B(n5295), .Y(n6253) );
   BF053  g843( .A1(n5463), .A2(n5460), .B1(n5228), .B2(
                           n6455), .Y(n5524) );
   EN210  g844( .A(n6252), .B(n6251), .Y(n6250) );
   IV110  g845( .A(n5524), .Y(n5523) );
   BF053  g846( .A1(n5420), .A2(n5419), .B1(n5239), .B2(
                           n5523), .Y(n5522) );
   EN210  g847( .A(n5991), .B(n6025), .Y(n6272) );
   BF003  g848( .A1(n5240), .A2(n5522), .B1(n5766), .B2(
                           n5312), .Y(n5521) );
   BF003  g849( .A1(n5875), .A2(n5276), .B1(n5992), .B2(
                           n5277), .Y(n6271) );
   BF053  g850( .A1(n5241), .A2(n5521), .B1(n6524), .B2(
                           n6523), .Y(n6476) );
   NA210  g851( .A(A_9_port), .B(B_12_port), .Y(n5917) );
   NA210  g853( .A(A_11_port), .B(B_10_port), .Y(n5918) );
   NA210  g854( .A(B_9_port), .B(A_12_port), .Y(n5919) );
   NA210  g855( .A(B_7_port), .B(A_14_port), .Y(n5660) );
   NA210  g856( .A(B_8_port), .B(A_14_port), .Y(n5661) );
   NA210  g857( .A(A_8_port), .B(B_14_port), .Y(n5662) );
   NA210  g858( .A(A_7_port), .B(B_15_port), .Y(n5663) );
   NA210  g859( .A(A_9_port), .B(B_13_port), .Y(n5664) );
   NA210  g860( .A(B_12_port), .B(A_10_port), .Y(n5665) );
   NA210  g861( .A(A_11_port), .B(B_11_port), .Y(n5666) );
   NA210  g862( .A(B_3_port), .B(A_10_port), .Y(n6416) );
   NO210  g863( .A(n5644), .B(n6418), .Y(n6417) );
   NA210  g864( .A(B_1_port), .B(A_6_port), .Y(n6419) );
   NO210  g865( .A(n6418), .B(n5557), .Y(n6420) );
   NA210  g866( .A(B_1_port), .B(A_8_port), .Y(n6421) );
   NO210  g867( .A(n6418), .B(n6423), .Y(n6422) );
   NA210  g868( .A(B_1_port), .B(A_10_port), .Y(n6424) );
   NO210  g869( .A(n6418), .B(n6176), .Y(n6425) );
   NA210  g870( .A(B_1_port), .B(A_12_port), .Y(n6177) );
   NA210  g871( .A(B_1_port), .B(A_13_port), .Y(n6178) );
   IV110  g872( .A(n6127), .Y(n6466) );
   NA210  g873( .A(B_5_port), .B(A_15_port), .Y(n5570) );
   IV110  g874( .A(n6183), .Y(n5880) );
   NO210  g875( .A(n6156), .B(n6157), .Y(n6160) );
   IV110  g876( .A(n5238), .Y(n5781) );
   AN210  g877( .A(n6159), .B(n6160), .Y(n5571) );
   IV110  g878( .A(n5656), .Y(n6303) );
   NO210  g879( .A(n5226), .B(n5652), .Y(n5572) );
   IV110  g880( .A(n5657), .Y(n6306) );
   NA210  g881( .A(B_4_port), .B(A_14_port), .Y(n5573) );
   BF003  g882( .A1(n6295), .A2(n6316), .B1(n5492), .B2(
                           n6317), .Y(n5541) );
   NA210  g883( .A(B_9_port), .B(A_6_port), .Y(n6077) );
   EN210  g884( .A(n5540), .B(n6365), .Y(n5544) );
   BF003  g885( .A1(n6294), .A2(n5889), .B1(n6363), .B2(
                           n6311), .Y(n5887) );
   EX210  g886( .A(n6364), .B(n5887), .Y(n5761) );
   BF053  g887( .A1(n5668), .A2(n5265), .B1(n6051), .B2(
                           n6050), .Y(n6326) );
   IV110  g888( .A(n6326), .Y(n6325) );
   BF053  g889( .A1(n6324), .A2(n5855), .B1(n6093), .B2(
                           n5800), .Y(n5920) );
   BF053  g890( .A1(n6086), .A2(n6325), .B1(n5856), .B2(
                           n5857), .Y(n6323) );
   IV110  g891( .A(n6323), .Y(n6322) );
   BF003  g892( .A1(n5436), .A2(n5594), .B1(n5480), .B2(
                           n5595), .Y(n5748) );
   NA210  g893( .A(A_4_port), .B(B_1_port), .Y(n5231) );
   EN210  g894( .A(n5747), .B(n5698), .Y(n6148) );
   NA210  g895( .A(A_2_port), .B(B_4_port), .Y(n5890) );
   EN210  g896( .A(n6264), .B(n6228), .Y(n6269) );
   NA210  g897( .A(n5455), .B(n6415), .Y(n5891) );
   BF003  g898( .A1(n5435), .A2(n5704), .B1(n5562), .B2(
                           n5706), .Y(n6268) );
   NO210  g899( .A(n6478), .B(n5232), .Y(n5894) );
   BF003  g900( .A1(n6395), .A2(n5280), .B1(n5994), .B2(
                           n5281), .Y(n5318) );
   NO210  g901( .A(n6175), .B(n5229), .Y(n5893) );
   BF053  g902( .A1(n6077), .A2(n6462), .B1(n6569), .B2(
                           n6570), .Y(n5604) );
   IV110  g903( .A(n5604), .Y(n5603) );
   BF053  g904( .A1(n6143), .A2(n6144), .B1(n6078), .B2(
                           n6465), .Y(n5602) );
   IV110  g905( .A(n5602), .Y(n5601) );
   BF053  g906( .A1(n6136), .A2(n6137), .B1(n6138), .B2(
                           n5739), .Y(n5600) );
   BF053  g907( .A1(n6079), .A2(n6556), .B1(n6557), .B2(
                           n6141), .Y(n6558) );
   BF003  g908( .A1(n5776), .A2(n6096), .B1(n5570), .B2(
                           n6097), .Y(n5755) );
   IV110  g909( .A(n6558), .Y(n6555) );
   EN210  g910( .A(n5624), .B(n5269), .Y(n6157) );
   BF053  g911( .A1(n6553), .A2(n6142), .B1(n6080), .B2(
                           n5514), .Y(n6554) );
   EN210  g912( .A(n6261), .B(n6260), .Y(n6259) );
   EN210  g913( .A(n6258), .B(n6257), .Y(n6256) );
   EN210  g914( .A(n5835), .B(n5838), .Y(n6255) );
   EN210  g915( .A(n6254), .B(n5839), .Y(n5838) );
   EN210  g916( .A(n5837), .B(n5836), .Y(n5835) );
   EX210  g917( .A(n5834), .B(n5833), .Y(n5832) );
   IV110  g918( .A(n6284), .Y(n6287) );
   EX210  g919( .A(n5831), .B(n5830), .Y(n5404) );
   BF053  g920( .A1(n5462), .A2(n5461), .B1(n5231), .B2(
                           n6449), .Y(n6288) );
   EX210  g921( .A(n5403), .B(n5402), .Y(n5401) );
   NO210  g922( .A(n6478), .B(n6184), .Y(n5837) );
   NO210  g923( .A(n6175), .B(n5982), .Y(n5836) );
   NA210  g924( .A(n5906), .B(n5905), .Y(n6254) );
   NA210  g925( .A(A_2_port), .B(B_12_port), .Y(n5839) );
   NA210  g926( .A(A_3_port), .B(B_11_port), .Y(n6185) );
   NA210  g927( .A(A_9_port), .B(B_10_port), .Y(n6433) );
   NA210  g928( .A(A_13_port), .B(B_7_port), .Y(n6434) );
   NA210  g929( .A(B_8_port), .B(A_12_port), .Y(n6435) );
   NA210  g930( .A(B_10_port), .B(A_10_port), .Y(n5475) );
   NA210  g931( .A(A_8_port), .B(B_12_port), .Y(n5476) );
   IV110  g932( .A(n5580), .Y(n5927) );
   NA210  g933( .A(A_2_port), .B(B_14_port), .Y(n6355) );
   IV110  g934( .A(n5925), .Y(n5583) );
   NA210  g935( .A(n6140), .B(n6139), .Y(n6356) );
   IV110  g936( .A(n5996), .Y(n5773) );
   NA210  g937( .A(n5924), .B(n5927), .Y(n6167) );
   IV110  g938( .A(n5577), .Y(n5775) );
   BF053  g939( .A1(n5974), .A2(n5975), .B1(n5973), .B2(
                           n5970), .Y(n6015) );
   IV110  g940( .A(n5578), .Y(n5774) );
   BF053  g941( .A1(n6448), .A2(n6413), .B1(n5227), .B2(
                           n6447), .Y(n6446) );
   IV110  g942( .A(n5979), .Y(n6196) );
   NA210  g943( .A(A_13_port), .B(B_10_port), .Y(n6092) );
   IV110  g944( .A(n5980), .Y(n5672) );
   IV110  g945( .A(n5985), .Y(n5678) );
   IV110  g946( .A(n5984), .Y(n5448) );
   BF056  g947( .A1(n5581), .A2(n6312), .B1(n5924), .B2(
                           n5536), .Y(n5342) );
   BF053  g948( .A1(n5542), .A2(n5541), .B1(n5492), .B2(
                           n6316), .Y(n5760) );
   BF053  g949( .A1(n5491), .A2(n6310), .B1(n5490), .B2(
                           n6313), .Y(n6311) );
   IV110  g950( .A(n6311), .Y(n5889) );
   NO210  g951( .A(n6366), .B(n5762), .Y(n5587) );
   EN210  g952( .A(n5857), .B(n5856), .Y(n5855) );
   EX2B0  g953( .A(n6274), .B(n5859), .Y(n5858) );
   EN210  g954( .A(n6277), .B(n6276), .Y(n6275) );
   EN210  g955( .A(n6280), .B(n6279), .Y(n6278) );
   EX210  g956( .A(n6283), .B(n6282), .Y(n6281) );
   EN210  g957( .A(n5327), .B(n5326), .Y(n5325) );
   EX210  g958( .A(n5329), .B(n5858), .Y(n5328) );
   EN2B0  g959( .A(n5462), .B(n5461), .Y(n5460) );
   EX2B0  g960( .A(n5332), .B(n5331), .Y(n5330) );
   EN210  g961( .A(n6414), .B(n5456), .Y(n5459) );
   BF053  g962( .A1(n6579), .A2(n6580), .B1(n5986), .B2(
                           n5284), .Y(n6226) );
   IV110  g963( .A(n6226), .Y(n5819) );
   BF053  g964( .A1(n5817), .A2(n5317), .B1(n5987), .B2(
                           n5283), .Y(n5818) );
   BF053  g965( .A1(n5815), .A2(n6273), .B1(n5988), .B2(
                           n6227), .Y(n5816) );
   IV110  g966( .A(n5816), .Y(n5814) );
   BF053  g967( .A1(n5989), .A2(n6230), .B1(n5812), .B2(
                           n6270), .Y(n5813) );
   IV110  g968( .A(n5813), .Y(n5811) );
   BF053  g969( .A1(n5990), .A2(n6233), .B1(n5991), .B2(
                           n6025), .Y(n5810) );
   IV110  g970( .A(n5810), .Y(n6024) );
   BF053  g971( .A1(n6272), .A2(n6271), .B1(n5992), .B2(
                           n5276), .Y(n6023) );
   NA210  g972( .A(B_3_port), .B(A_9_port), .Y(n6494) );
   NA210  g973( .A(B_4_port), .B(A_8_port), .Y(n6495) );
   NA210  g974( .A(B_5_port), .B(A_7_port), .Y(n6496) );
   NA210  g975( .A(B_6_port), .B(A_6_port), .Y(n6497) );
   NA210  g976( .A(A_4_port), .B(B_8_port), .Y(n6498) );
   NO210  g977( .A(n6478), .B(n5550), .Y(n5721) );
   NO210  g978( .A(n6175), .B(n6492), .Y(n5720) );
   NA210  g979( .A(n6252), .B(n6251), .Y(n5724) );
   NA210  g980( .A(A_2_port), .B(B_10_port), .Y(n5723) );
   NA210  g981( .A(A_3_port), .B(B_9_port), .Y(n5551) );
   EN210  g982( .A(n5630), .B(n6592), .Y(n5224) );
   BF001  g983( .A1(n6241), .B1(n5533), .B2(n6240), .Y(
                           n6239) );
   BF003  g984( .A1(n5633), .A2(n5632), .B1(n5635), .B2(
                           n5634), .Y(n5631) );
   BF006  g985( .A1(n6238), .A2(n6381), .B1(n6237), .B2(
                           n5944), .Y(n6236) );
   NO210  g986( .A(n5539), .B(n5538), .Y(n5537) );
   NO210  g987( .A(n5536), .B(n5535), .Y(n5534) );
   NA210  g988( .A(n5533), .B(n5532), .Y(n5531) );
   NO210  g989( .A(n6478), .B(n6477), .Y(PRODUCT_0_port) );
   BF001  g990( .A1(n6385), .B1(n6384), .B2(n6383), .Y(
                           PRODUCT_18_port) );
   NO210  g991( .A(n5644), .B(n5226), .Y(n5643) );
   IV110  g992( .A(n5988), .Y(n5871) );
   BF053  g993( .A1(n5486), .A2(n6314), .B1(n5485), .B2(
                           n6319), .Y(n6315) );
   IV110  g994( .A(n5995), .Y(n5953) );
   IV110  g995( .A(n6315), .Y(n6313) );
   IV110  g996( .A(n6433), .Y(n5441) );
   IV110  g997( .A(n6432), .Y(n5442) );
   IV110  g998( .A(n6430), .Y(n5443) );
   IV110  g999( .A(n6429), .Y(n5444) );
   IV110  g1000( .A(n6428), .Y(n5870) );
   IV110  g1001( .A(n6427), .Y(n6394) );
   BF053  g1002( .A1(n5476), .A2(n6545), .B1(n5695), .B2(
                           n5744), .Y(n5696) );
   IV110  g1003( .A(n5696), .Y(n5694) );
   BF053  g1004( .A1(n5478), .A2(n5692), .B1(n5477), .B2(
                           n6548), .Y(n5693) );
   IV110  g1005( .A(n5693), .Y(n5691) );
   BF053  g1006( .A1(n5479), .A2(n5592), .B1(n5746), .B2(
                           n5745), .Y(n5690) );
   IV110  g1007( .A(n5690), .Y(n5274) );
   IV110  g1008( .A(n5641), .Y(n6201) );
   BF053  g1009( .A1(n5480), .A2(n5594), .B1(n5749), .B2(
                           n5748), .Y(n5273) );
   IV110  g1010( .A(n5645), .Y(n5676) );
   IV110  g1011( .A(n5273), .Y(n5272) );
   EN210  g1012( .A(n6330), .B(n5899), .Y(n5898) );
   EN210  g1013( .A(n5897), .B(n5896), .Y(n5895) );
   EN210  g1014( .A(n5894), .B(n5893), .Y(n5892) );
   EN210  g1015( .A(n5891), .B(n5890), .Y(n5464) );
   NO210  g1016( .A(n6175), .B(n5226), .Y(n6415) );
   EX210  g1017( .A(n5460), .B(n5463), .Y(PRODUCT_5_port) );
   NA210  g1018( .A(n6409), .B(n6408), .Y(n5458) );
   NA210  g1019( .A(A_2_port), .B(B_3_port), .Y(n5457) );
   EN210  g1020( .A(n5744), .B(n5695), .Y(n5749) );
   NA210  g1021( .A(A_3_port), .B(B_2_port), .Y(n5230) );
   IV110  g1022( .A(n5600), .Y(n6117) );
   IV110  g1023( .A(n6499), .Y(n5246) );
   IV110  g1024( .A(n6085), .Y(n5247) );
   IV110  g1025( .A(n6084), .Y(n5248) );
   IV110  g1026( .A(n5568), .Y(n5872) );
   EN210  g1027( .A(n6259), .B(n5519), .Y(n5305) );
   BF003  g1028( .A1(n5676), .A2(n5429), .B1(n5645), .B2(
                           n5939), .Y(n5428) );
   BF003  g1029( .A1(n5675), .A2(n5430), .B1(n6072), .B2(
                           n5427), .Y(n6245) );
   EN210  g1030( .A(n5829), .B(n6285), .Y(n6246) );
   BF003  g1031( .A1(n5674), .A2(n5868), .B1(n6490), .B2(
                           n5867), .Y(n5962) );
   IV110  g1032( .A(n5591), .Y(n6548) );
   IV110  g1033( .A(B_0_port), .Y(n6477) );
   BF053  g1034( .A1(n6432), .A2(n5811), .B1(n6546), .B2(
                           n5320), .Y(n6547) );
   IV110  g1035( .A(B_8_port), .Y(n5642) );
   IV110  g1036( .A(n6547), .Y(n6545) );
   IV110  g1037( .A(A_9_port), .Y(n6423) );
   BF053  g1038( .A1(n6433), .A2(n5814), .B1(n6543), .B2(
                           n5323), .Y(n6544) );
   IV110  g1039( .A(A_7_port), .Y(n5557) );
   IV110  g1040( .A(n6544), .Y(n6542) );
   IV110  g1041( .A(A_5_port), .Y(n5644) );
   IV110  g1042( .A(n6129), .Y(n6128) );
   BF053  g1043( .A1(n5908), .A2(n5909), .B1(n5907), .B2(
                           n5904), .Y(n6127) );
   BF053  g1044( .A1(n5983), .A2(n5718), .B1(n5719), .B2(
                           n6340), .Y(n6126) );
   IV110  g1045( .A(n6126), .Y(n5717) );
   BF053  g1046( .A1(n5978), .A2(n6468), .B1(n5715), .B2(
                           n6347), .Y(n5716) );
   BF053  g1047( .A1(n5563), .A2(n5707), .B1(n6265), .B2(
                           n6266), .Y(n5279) );
   IV110  g1048( .A(n5279), .Y(n5278) );
   BF053  g1049( .A1(n5564), .A2(n6116), .B1(n5848), .B2(
                           n5849), .Y(n5277) );
   IV110  g1050( .A(n5277), .Y(n5276) );
   BF053  g1051( .A1(n5565), .A2(n6234), .B1(n5566), .B2(
                           n6235), .Y(n5275) );
   EN210  g1052( .A(n5841), .B(n5680), .Y(n5846) );
   EN210  g1053( .A(n5306), .B(n5290), .Y(n5311) );
   EN210  g1054( .A(n6247), .B(n5861), .Y(n5831) );
   EN210  g1055( .A(n5394), .B(n5502), .Y(n5400) );
   BF003  g1056( .A1(n5356), .A2(n5498), .B1(n5553), .B2(
                           n5495), .Y(n5399) );
   EN210  g1057( .A(n6488), .B(n6487), .Y(n6486) );
   EX210  g1058( .A(n5542), .B(n5541), .Y(n5540) );
   EN210  g1059( .A(n5545), .B(n5544), .Y(n5543) );
   EN210  g1060( .A(n5548), .B(n5547), .Y(n5546) );
   EX2B0  g1061( .A(n5336), .B(n5335), .Y(n5549) );
   IV110  g1062( .A(n6013), .Y(n5585) );
   BF053  g1063( .A1(n5661), .A2(n5803), .B1(n5801), .B2(
                           n6049), .Y(n5802) );
   IV110  g1064( .A(n6015), .Y(n6447) );
   IV110  g1065( .A(n5802), .Y(n5800) );
   IV110  g1066( .A(n5231), .Y(n5882) );
   IV110  g1067( .A(n6450), .Y(n5496) );
   IV110  g1068( .A(n6452), .Y(n6454) );
   IV110  g1069( .A(n5228), .Y(n5884) );
   IV110  g1070( .A(n5553), .Y(n5356) );
   IV110  g1071( .A(n5503), .Y(n5934) );
   EN210  g1072( .A(n6270), .B(n5812), .Y(n5316) );
   BF003  g1073( .A1(n5242), .A2(n6476), .B1(n6057), .B2(
                           n5730), .Y(n6475) );
   EN210  g1074( .A(n5847), .B(n6231), .Y(n6266) );
   BF053  g1075( .A1(n5418), .A2(n5417), .B1(n5243), .B2(
                           n6475), .Y(n6474) );
   BF003  g1076( .A1(n5874), .A2(n5707), .B1(n5563), .B2(
                           n5709), .Y(n6265) );
   BF003  g1077( .A1(n5873), .A2(n5278), .B1(n5993), .B2(
                           n5279), .Y(n5315) );
   BF003  g1078( .A1(n5872), .A2(n6123), .B1(n5568), .B2(
                           n6124), .Y(n6228) );
   BF003  g1079( .A1(n5871), .A2(n6227), .B1(n5988), .B2(
                           n6229), .Y(n5815) );
   BF003  g1080( .A1(n5870), .A2(n6020), .B1(n6428), .B2(
                           n6021), .Y(n5324) );
   BF003  g1081( .A1(n5444), .A2(n6022), .B1(n6429), .B2(
                           n6023), .Y(n5321) );
   NA210  g1082( .A(n5920), .B(n6281), .Y(n5340) );
   NO210  g1083( .A(n5546), .B(n5340), .Y(n5921) );
   NA210  g1084( .A(n5549), .B(n5921), .Y(n5922) );
   OR210  g1085( .A(n5326), .B(n5327), .Y(n5923) );
   NA210  g1086( .A(n5328), .B(n5571), .Y(n5924) );
   NO210  g1087( .A(n5325), .B(n6515), .Y(n5535) );
   NA410  g1088( .A(n5533), .B(n5926), .C(n5927), .D(n5928), 
                           .Y(n5925) );
   BF056  g1089( .A1(n6362), .A2(n6361), .B1(n6360), .B2(
                           n5539), .Y(n5929) );
   NA210  g1090( .A(A_15_port), .B(B_14_port), .Y(n6363) );
   NA210  g1091( .A(A_14_port), .B(B_15_port), .Y(n6364) );
   NA210  g1092( .A(A_7_port), .B(B_11_port), .Y(n5993) );
   NA210  g1093( .A(A_9_port), .B(B_9_port), .Y(n5994) );
   NA210  g1094( .A(B_7_port), .B(A_12_port), .Y(n5995) );
   NO210  g1095( .A(n6176), .B(n5642), .Y(n6426) );
   NA210  g1096( .A(B_9_port), .B(A_10_port), .Y(n6427) );
   NA210  g1097( .A(A_8_port), .B(B_11_port), .Y(n6428) );
   NA210  g1098( .A(A_6_port), .B(B_13_port), .Y(n6429) );
   NA210  g1099( .A(A_5_port), .B(B_14_port), .Y(n6430) );
   NA210  g1100( .A(A_4_port), .B(B_15_port), .Y(n6431) );
   NA210  g1101( .A(A_7_port), .B(B_12_port), .Y(n6432) );
   IV110  g1102( .A(n5658), .Y(n5358) );
   NO210  g1103( .A(n5226), .B(n5655), .Y(n5574) );
   IV110  g1104( .A(n5659), .Y(n5780) );
   IV110  g1105( .A(n6076), .Y(n5249) );
   IV110  g1106( .A(n6082), .Y(n5250) );
   BF002  g1107( .A1(n5535), .B1(n5533), .B2(n6240), .B3(
                           n6528), .Y(n5581) );
   BF002  g1108( .A1(n5585), .B1(n6240), .B2(n5583), .B3(
                           n5584), .Y(n5582) );
   BF052  g1109( .A1(n5588), .B1(n6382), .B2(n5416), .B3(
                           n5587), .Y(n5586) );
   IV110  g1110( .A(n6514), .Y(n5352) );
   BF001  g1111( .A1(n5586), .B1(n5929), .B2(n5584), .Y(
                           n5589) );
   BF053  g1112( .A1(n6320), .A2(n5852), .B1(n6092), .B2(
                           n5382), .Y(n6321) );
   IV110  g1113( .A(n5863), .Y(n6398) );
   IV110  g1114( .A(n6321), .Y(n6538) );
   IV110  g1115( .A(n6489), .Y(n6198) );
   BF053  g1116( .A1(n5854), .A2(n5853), .B1(n6091), .B2(
                           n5380), .Y(n6537) );
   IV110  g1117( .A(n6490), .Y(n5674) );
   IV110  g1118( .A(n6537), .Y(n6536) );
   IV110  g1119( .A(n5869), .Y(n5530) );
   BF053  g1120( .A1(n6534), .A2(n6055), .B1(n6090), .B2(
                           n5377), .Y(n6535) );
   IV110  g1121( .A(n6491), .Y(n5445) );
   EN210  g1122( .A(n6273), .B(n5815), .Y(n5319) );
   NA210  g1123( .A(A_3_port), .B(B_4_port), .Y(n5233) );
   EN210  g1124( .A(n5323), .B(n6543), .Y(n5743) );
   BF003  g1125( .A1(n6394), .A2(n6018), .B1(n6427), .B2(
                           n6019), .Y(n5742) );
   BF003  g1126( .A1(n6393), .A2(n5596), .B1(n5481), .B2(
                           n5597), .Y(n6147) );
   IV110  g1127( .A(n6551), .Y(n6549) );
   BF053  g1128( .A1(n6503), .A2(n5605), .B1(n5412), .B2(
                           n5411), .Y(n6125) );
   BF053  g1129( .A1(n6085), .A2(n6552), .B1(n5408), .B2(
                           n5409), .Y(n6124) );
   IV110  g1130( .A(n6124), .Y(n6123) );
   BF053  g1131( .A1(n6499), .A2(n6555), .B1(n5405), .B2(
                           n5406), .Y(n6122) );
   BF003  g1132( .A1(n6417), .A2(n6288), .B1(n6290), .B2(
                           n5398), .Y(n6289) );
   EX210  g1133( .A(n5400), .B(n5399), .Y(n5398) );
   BF053  g1134( .A1(n5314), .A2(n5313), .B1(n6419), .B2(
                           n6289), .Y(n6291) );
   EN210  g1135( .A(n5397), .B(n5396), .Y(n5395) );
   BF003  g1136( .A1(n6293), .A2(n5401), .B1(n6420), .B2(
                           n6291), .Y(n6292) );
   BF053  g1137( .A1(n5731), .A2(n5732), .B1(n6421), .B2(
                           n6292), .Y(n6405) );
   BF003  g1138( .A1(n6301), .A2(n5523), .B1(n5239), .B2(
                           n5524), .Y(n5420) );
   BF003  g1139( .A1(n6403), .A2(n5404), .B1(n6422), .B2(
                           n6405), .Y(n6404) );
   EX210  g1140( .A(n5240), .B(n5522), .Y(n5766) );
   BF053  g1141( .A1(n5735), .A2(n5734), .B1(n6424), .B2(
                           n6404), .Y(n6402) );
   NA210  g1142( .A(A_6_port), .B(B_14_port), .Y(n5477) );
   NA210  g1143( .A(A_5_port), .B(B_15_port), .Y(n5478) );
   NA210  g1144( .A(A_7_port), .B(B_13_port), .Y(n5479) );
   NA210  g1145( .A(A_9_port), .B(B_11_port), .Y(n5480) );
   NA210  g1146( .A(A_11_port), .B(B_9_port), .Y(n5481) );
   NA210  g1147( .A(B_13_port), .B(A_12_port), .Y(n6438) );
   NA210  g1148( .A(A_11_port), .B(B_14_port), .Y(n6439) );
   NA210  g1149( .A(A_10_port), .B(B_15_port), .Y(n6440) );
   NA210  g1150( .A(A_15_port), .B(B_11_port), .Y(n6441) );
   AN210  g1151( .A(B_12_port), .B(A_14_port), .Y(n6442) );
   NA410  g1152( .A(n6368), .B(n5941), .C(n5415), .D(n6237), 
                           .Y(n5588) );
   IV110  g1153( .A(n5917), .Y(n6388) );
   BF056  g1154( .A1(n5589), .A2(n5582), .B1(n5888), .B2(
                           n5587), .Y(n5423) );
   IV110  g1155( .A(n5915), .Y(n6389) );
   BF053  g1156( .A1(n6364), .A2(n5887), .B1(n6363), .B2(
                           n5889), .Y(n6009) );
   IV110  g1157( .A(n5914), .Y(n6390) );
   NA410  g1158( .A(n6369), .B(n5769), .C(n5415), .D(n6237), 
                           .Y(n6010) );
   IV110  g1159( .A(n5913), .Y(n6391) );
   BF001  g1160( .A1(n6004), .B1(n6385), .B2(n6011), .Y(
                           n6168) );
   IV110  g1161( .A(n5660), .Y(n5951) );
   EN210  g1162( .A(n5750), .B(n5334), .Y(n5333) );
   EN210  g1163( .A(n5458), .B(n5457), .Y(n5456) );
   EX210  g1164( .A(n5753), .B(n5752), .Y(n5751) );
   EN210  g1165( .A(n5455), .B(n6415), .Y(n6414) );
   EN210  g1166( .A(n6407), .B(n6410), .Y(n6413) );
   EN210  g1167( .A(n6412), .B(n6411), .Y(n6410) );
   EN210  g1168( .A(n6409), .B(n6408), .Y(n6407) );
   EN210  g1169( .A(n5970), .B(n5973), .Y(n6406) );
   EN210  g1170( .A(n5975), .B(n5974), .Y(n5973) );
   NA210  g1171( .A(n5894), .B(n5893), .Y(n5897) );
   NA210  g1172( .A(B_6_port), .B(A_10_port), .Y(n6084) );
   NA210  g1173( .A(A_6_port), .B(B_10_port), .Y(n6085) );
   NA210  g1174( .A(A_4_port), .B(B_12_port), .Y(n6499) );
   NA210  g1175( .A(A_1_port), .B(B_15_port), .Y(n6358) );
   NA210  g1176( .A(A_3_port), .B(B_13_port), .Y(n6500) );
   NA210  g1177( .A(A_5_port), .B(B_11_port), .Y(n6501) );
   NA210  g1178( .A(A_7_port), .B(B_9_port), .Y(n6502) );
   NA210  g1179( .A(A_8_port), .B(B_8_port), .Y(n6503) );
   NA210  g1180( .A(A_9_port), .B(B_7_port), .Y(n6504) );
   NA210  g1181( .A(B_5_port), .B(A_11_port), .Y(n6505) );
   NO210  g1182( .A(n6382), .B(n6381), .Y(n6380) );
   NA210  g1183( .A(A_3_port), .B(B_6_port), .Y(n5645) );
   NO210  g1184( .A(n6478), .B(n5646), .Y(n5386) );
   EN210  g1185( .A(n6584), .B(n6219), .Y(n5620) );
   NO210  g1186( .A(n6175), .B(n5642), .Y(n5385) );
   BF003  g1187( .A1(n6387), .A2(n5697), .B1(n5918), .B2(
                           n5699), .Y(n6224) );
   NA210  g1188( .A(n6337), .B(n6336), .Y(n5389) );
   EN210  g1189( .A(n6587), .B(n6224), .Y(n5623) );
   NA210  g1190( .A(A_2_port), .B(B_7_port), .Y(n5388) );
   BF003  g1191( .A1(n6386), .A2(n6106), .B1(n5919), .B2(
                           n6107), .Y(n5622) );
   BF003  g1192( .A1(n5247), .A2(n6552), .B1(n6085), .B2(
                           n6554), .Y(n5408) );
   BF003  g1193( .A1(n5246), .A2(n6555), .B1(n6499), .B2(
                           n6558), .Y(n5405) );
   BF003  g1194( .A1(n5245), .A2(n6117), .B1(n6500), .B2(
                           n5600), .Y(n6118) );
   EN210  g1195( .A(n6357), .B(n6118), .Y(n5406) );
   BF003  g1196( .A1(n6205), .A2(n5601), .B1(n6501), .B2(
                           n5602), .Y(n5708) );
   EN210  g1197( .A(n6359), .B(n5708), .Y(n5409) );
   BF003  g1198( .A1(n6204), .A2(n5603), .B1(n6502), .B2(
                           n5604), .Y(n5705) );
   EN210  g1199( .A(n5407), .B(n5705), .Y(n5412) );
   BF003  g1200( .A1(n6203), .A2(n5605), .B1(n6503), .B2(
                           n5607), .Y(n5411) );
   BF003  g1201( .A1(n6202), .A2(n5608), .B1(n6504), .B2(
                           n5609), .Y(n5702) );
   IV110  g1202( .A(n6068), .Y(n5363) );
   BF053  g1203( .A1(n6434), .A2(n6016), .B1(n6150), .B2(
                           n6151), .Y(n5271) );
   IV110  g1204( .A(n6071), .Y(n5446) );
   IV110  g1205( .A(n5271), .Y(n5270) );
   IV110  g1206( .A(n6075), .Y(n5784) );
   IV110  g1207( .A(n6493), .Y(n5450) );
   IV110  g1208( .A(n5551), .Y(n5453) );
   IV110  g1209( .A(n5559), .Y(n5355) );
   IV110  g1210( .A(n5983), .Y(n5881) );
   IV110  g1211( .A(n6178), .Y(n6304) );
   BF053  g1212( .A1(n6263), .A2(n5305), .B1(n6182), .B2(
                           n6135), .Y(n5286) );
   IV110  g1213( .A(n5286), .Y(n5285) );
   BF053  g1214( .A1(n5519), .A2(n6259), .B1(n5237), .B2(
                           n6133), .Y(n5520) );
   IV110  g1215( .A(n5520), .Y(n5518) );
   BF053  g1216( .A1(n6261), .A2(n6260), .B1(n5236), .B2(
                           n6130), .Y(n5517) );
   IV110  g1217( .A(n5517), .Y(n5516) );
   BF003  g1218( .A1(n5949), .A2(n5807), .B1(n5662), .B2(
                           n5809), .Y(n6328) );
   BF053  g1219( .A1(n6257), .A2(n6258), .B1(n6183), .B2(
                           n5717), .Y(n5515) );
   EN210  g1220( .A(n5663), .B(n6328), .Y(n5629) );
   IV110  g1221( .A(n5515), .Y(n5514) );
   EN210  g1222( .A(n5726), .B(n6040), .Y(n5466) );
   BF003  g1223( .A1(n5673), .A2(n5961), .B1(n6497), .B2(
                           n5963), .Y(n5465) );
   BF003  g1224( .A1(n5672), .A2(n6042), .B1(n5980), .B2(
                           n6043), .Y(n6559) );
   BF003  g1225( .A1(n5671), .A2(n6135), .B1(n6182), .B2(
                           n6560), .Y(n6263) );
   BF003  g1226( .A1(n5670), .A2(n6462), .B1(n6077), .B2(
                           n6464), .Y(n6569) );
   EX2B0  g1227( .A(n5422), .B(n5421), .Y(PRODUCT_14_port) );
   EX210  g1228( .A(n5424), .B(n5423), .Y(PRODUCT_30_port) );
   EX2B0  g1229( .A(n6520), .B(n6519), .Y(PRODUCT_4_port) );
   EX2B0  g1230( .A(n6522), .B(n6521), .Y(PRODUCT_12_port) );
   EX2B0  g1231( .A(n6170), .B(n6171), .Y(PRODUCT_1_port) );
   IV110  g1232( .A(B_6_port), .Y(n5232) );
   IV110  g1233( .A(B_1_port), .Y(n6418) );
   IV110  g1234( .A(B_4_port), .Y(n5226) );
   IV110  g1235( .A(B_7_port), .Y(n5234) );
   IV110  g1236( .A(A_1_port), .Y(n6175) );
   BF053  g1237( .A1(n6517), .A2(n6100), .B1(n5334), .B2(
                           n5750), .Y(n6099) );
   IV110  g1238( .A(n6099), .Y(n6098) );
   BF053  g1239( .A1(n5331), .A2(n5332), .B1(n6518), .B2(
                           n6098), .Y(n6097) );
   IV110  g1240( .A(n6097), .Y(n6096) );
   BF053  g1241( .A1(n5755), .A2(n5756), .B1(n5570), .B2(
                           n6096), .Y(n5758) );
   IV110  g1242( .A(n5275), .Y(n6233) );
   BF053  g1243( .A1(n6231), .A2(n5847), .B1(n5567), .B2(
                           n6121), .Y(n6232) );
   IV110  g1244( .A(n6232), .Y(n6230) );
   BF053  g1245( .A1(n5568), .A2(n6123), .B1(n6228), .B2(
                           n6264), .Y(n6229) );
   IV110  g1246( .A(n6229), .Y(n6227) );
   OR210  g1247( .A(n5969), .B(n5968), .Y(n5975) );
   NA210  g1248( .A(B_1_port), .B(A_2_port), .Y(n5974) );
   NA210  g1249( .A(B_0_port), .B(A_4_port), .Y(n5225) );
   NO210  g1250( .A(n6478), .B(n5226), .Y(n6409) );
   NO210  g1251( .A(n6175), .B(n6173), .Y(n6408) );
   EX210  g1252( .A(n5338), .B(n6486), .Y(n5337) );
   EN210  g1253( .A(n5340), .B(n5546), .Y(n5339) );
   EX210  g1254( .A(n6380), .B(n5341), .Y(PRODUCT_28_port) );
   EX210  g1255( .A(n5537), .B(n5342), .Y(PRODUCT_25_port) );
   EX2B0  g1256( .A(n6406), .B(n5343), .Y(PRODUCT_3_port) );
   NA210  g1257( .A(B_3_port), .B(A_8_port), .Y(n6074) );
   NA210  g1258( .A(B_4_port), .B(A_7_port), .Y(n6075) );
   NA210  g1259( .A(B_5_port), .B(A_6_port), .Y(n6489) );
   NA210  g1260( .A(A_5_port), .B(B_6_port), .Y(n6490) );
   NA210  g1261( .A(A_4_port), .B(B_7_port), .Y(n6491) );
   EN210  g1262( .A(n5729), .B(n6045), .Y(n5469) );
   BF003  g1263( .A1(n5786), .A2(n5934), .B1(n5233), .B2(
                           n5503), .Y(n5935) );
   BF003  g1264( .A1(n5785), .A2(n5936), .B1(n5640), .B2(
                           n5933), .Y(n5821) );
   EN210  g1265( .A(n6338), .B(n6371), .Y(n5822) );
   EX2B0  g1266( .A(n5938), .B(n5643), .Y(n5432) );
   IV110  g1267( .A(n5798), .Y(n5796) );
   BF053  g1268( .A1(n5795), .A2(n6061), .B1(n6005), .B2(
                           n6212), .Y(n5489) );
   BF053  g1269( .A1(n6062), .A2(n6063), .B1(n6436), .B2(
                           n6210), .Y(n5794) );
   IV110  g1270( .A(n5794), .Y(n5793) );
   BF053  g1271( .A1(n6437), .A2(n6207), .B1(n5791), .B2(
                           n6058), .Y(n5792) );
   BF053  g1272( .A1(n6059), .A2(n6060), .B1(n6438), .B2(
                           n5799), .Y(n5790) );
   IV110  g1273( .A(n5567), .Y(n5878) );
   IV110  g1274( .A(n5790), .Y(n5374) );
   IV110  g1275( .A(n6120), .Y(n6234) );
   BF053  g1276( .A1(n6440), .A2(n5372), .B1(n6439), .B2(
                           n5796), .Y(n5373) );
   BF053  g1277( .A1(n6578), .A2(n6350), .B1(n5658), .B2(
                           n5289), .Y(n6032) );
   IV110  g1278( .A(n6032), .Y(n6031) );
   BF053  g1279( .A1(n6029), .A2(n6574), .B1(n5659), .B2(
                           n5287), .Y(n6030) );
   IV110  g1280( .A(n6030), .Y(n6028) );
   BF053  g1281( .A1(n6576), .A2(n6575), .B1(n6083), .B2(
                           n6459), .Y(n6027) );
   IV110  g1282( .A(n6027), .Y(n6026) );
   BF003  g1283( .A1(n6186), .A2(n5800), .B1(n6093), .B2(
                           n5802), .Y(n6324) );
   BF053  g1284( .A1(n6573), .A2(n6572), .B1(n6082), .B2(
                           n5518), .Y(n5609) );
   EX210  g1285( .A(n5855), .B(n6324), .Y(n6274) );
   IV110  g1286( .A(n5609), .Y(n5608) );
   EN210  g1287( .A(n6138), .B(n5739), .Y(n6141) );
   EN210  g1288( .A(n6140), .B(n6139), .Y(n6138) );
   EN210  g1289( .A(n6137), .B(n6136), .Y(n5739) );
   EX210  g1290( .A(n5738), .B(n5737), .Y(n5736) );
   EX210  g1291( .A(n5735), .B(n5734), .Y(n5733) );
   EX210  g1292( .A(n5732), .B(n5731), .Y(n5730) );
   BF053  g1293( .A1(n5830), .A2(n5831), .B1(n5558), .B2(
                           n6376), .Y(n5433) );
   EX210  g1294( .A(n5314), .B(n5313), .Y(n5312) );
   BF053  g1295( .A1(n5861), .A2(n6247), .B1(n6068), .B2(
                           n5860), .Y(n5434) );
   EN210  g1296( .A(n5311), .B(n5310), .Y(n5309) );
   NA210  g1297( .A(n5631), .B(n5997), .Y(n6384) );
   NA210  g1298( .A(n6000), .B(n6589), .Y(n5630) );
   NO210  g1299( .A(n6383), .B(n6384), .Y(n6385) );
   NO210  g1300( .A(n6592), .B(n5630), .Y(n6001) );
   NA210  g1301( .A(n5221), .B(n6001), .Y(n6002) );
   NA210  g1302( .A(n5636), .B(n5637), .Y(n6003) );
   NO210  g1303( .A(n5224), .B(n6003), .Y(n6004) );
   NA210  g1304( .A(A_15_port), .B(B_10_port), .Y(n6005) );
   NA210  g1305( .A(B_11_port), .B(A_14_port), .Y(n6436) );
   NA210  g1306( .A(A_13_port), .B(B_12_port), .Y(n6437) );
   NA210  g1307( .A(A_13_port), .B(B_11_port), .Y(n6512) );
   IV110  g1308( .A(n6179), .Y(n6307) );
   NA210  g1309( .A(B_10_port), .B(A_14_port), .Y(n6513) );
   IV110  g1310( .A(n6180), .Y(n5359) );
   NA210  g1311( .A(A_15_port), .B(B_9_port), .Y(n6514) );
   IV110  g1312( .A(n6181), .Y(n5789) );
   NA210  g1313( .A(n5859), .B(n6274), .Y(n5327) );
   IV110  g1314( .A(n6182), .Y(n5671) );
   IV110  g1315( .A(n5237), .Y(n5677) );
   IV110  g1316( .A(n5236), .Y(n5447) );
   IV110  g1317( .A(n6513), .Y(n5353) );
   EX2B0  g1318( .A(n6008), .B(n6007), .Y(n6006) );
   IV110  g1319( .A(n6512), .Y(n5354) );
   EX210  g1320( .A(n6009), .B(n6006), .Y(n5424) );
   IV110  g1321( .A(n6511), .Y(n5770) );
   BF052  g1322( .A1(n6010), .B1(n6382), .B2(n5922), .B3(
                           n5945), .Y(n6238) );
   IV110  g1323( .A(n6510), .Y(n5771) );
   NA210  g1324( .A(n6012), .B(n6011), .Y(n6525) );
   IV110  g1325( .A(n6095), .Y(n5772) );
   NA210  g1326( .A(n6161), .B(n5579), .Y(n5509) );
   IV110  g1327( .A(n6494), .Y(n5361) );
   IV110  g1328( .A(n6495), .Y(n5783) );
   IV110  g1329( .A(n6496), .Y(n6197) );
   IV110  g1330( .A(n6497), .Y(n5673) );
   IV110  g1331( .A(n5552), .Y(n5679) );
   NA210  g1332( .A(n5493), .B(n5543), .Y(n6237) );
   BF053  g1333( .A1(n6283), .A2(n6282), .B1(n6514), .B2(
                           n6322), .Y(n5548) );
   NO210  g1334( .A(n5494), .B(n5337), .Y(n5945) );
   NO210  g1335( .A(n5921), .B(n5549), .Y(n5942) );
   NA210  g1336( .A(n5923), .B(n5339), .Y(n5926) );
   IV110  g1337( .A(n6122), .Y(n6121) );
   EX2B0  g1338( .A(n5330), .B(n5684), .Y(n5220) );
   BF051  g1339( .A1(n6356), .B1(n6358), .B2(n6354), .Y(
                           n6120) );
   BF003  g1340( .A1(n5773), .A2(n5682), .B1(n5996), .B2(
                           n5683), .Y(n5263) );
   BF053  g1341( .A1(n6500), .A2(n6117), .B1(n6118), .B2(
                           n6357), .Y(n6119) );
   EX210  g1342( .A(n6589), .B(n6000), .Y(n5636) );
   IV110  g1343( .A(n6119), .Y(n6116) );
   EN210  g1344( .A(n6163), .B(n5263), .Y(n5635) );
   BF053  g1345( .A1(n5708), .A2(n6359), .B1(n6501), .B2(
                           n5601), .Y(n5709) );
   BF003  g1346( .A1(n5772), .A2(n6105), .B1(n6095), .B2(
                           n6530), .Y(n5797) );
   EN210  g1347( .A(n5906), .B(n5905), .Y(n5904) );
   BF053  g1348( .A1(n6397), .A2(n5301), .B1(n6075), .B2(
                           n6398), .Y(n6399) );
   EN210  g1349( .A(n5903), .B(n5902), .Y(n5901) );
   IV110  g1350( .A(n6399), .Y(n6396) );
   EX210  g1351( .A(n5900), .B(n5474), .Y(n5473) );
   BF053  g1352( .A1(n6489), .A2(n5866), .B1(n5302), .B2(
                           n5303), .Y(n5965) );
   EX210  g1353( .A(n5472), .B(n5471), .Y(n5470) );
   IV110  g1354( .A(n5965), .Y(n5964) );
   EN210  g1355( .A(n5469), .B(n5468), .Y(n5467) );
   BF053  g1356( .A1(n6490), .A2(n5868), .B1(n5962), .B2(
                           n5298), .Y(n5963) );
   EN210  g1357( .A(n5401), .B(n6293), .Y(n6523) );
   BF053  g1358( .A1(n5902), .A2(n5903), .B1(n6074), .B2(
                           n5862), .Y(n6401) );
   EN210  g1359( .A(n5241), .B(n5521), .Y(n6524) );
   IV110  g1360( .A(n6401), .Y(n6400) );
   EX2B0  g1361( .A(n5242), .B(n6476), .Y(n6057) );
   EN2B0  g1362( .A(n5243), .B(n6475), .Y(n5417) );
   EN210  g1363( .A(n5404), .B(n6403), .Y(n5418) );
   EX210  g1364( .A(n5244), .B(n6474), .Y(n5764) );
   EN2B0  g1365( .A(n5650), .B(n6473), .Y(n6521) );
   EN2B0  g1366( .A(n5832), .B(n5611), .Y(n6522) );
   NA210  g1367( .A(A_13_port), .B(B_13_port), .Y(n6443) );
   NA210  g1368( .A(A_12_port), .B(B_14_port), .Y(n6444) );
   NA210  g1369( .A(A_11_port), .B(B_15_port), .Y(n6445) );
   NA210  g1370( .A(A_13_port), .B(B_14_port), .Y(n5485) );
   NA210  g1371( .A(A_12_port), .B(B_15_port), .Y(n5486) );
   BF053  g1372( .A1(n5891), .A2(n5890), .B1(n5892), .B2(
                           n5464), .Y(n5503) );
   BF003  g1373( .A1(n5554), .A2(n5500), .B1(n5930), .B2(
                           n5470), .Y(n5504) );
   BF053  g1374( .A1(n5471), .A2(n5472), .B1(n5649), .B2(
                           n5501), .Y(n5931) );
   BF053  g1375( .A1(n5896), .A2(n5897), .B1(n5898), .B2(
                           n5895), .Y(n5932) );
   BF053  g1376( .A1(n5935), .A2(n6331), .B1(n5233), .B2(
                           n5934), .Y(n5933) );
   IV110  g1377( .A(n5669), .Y(n6193) );
   IV110  g1378( .A(n5668), .Y(n6194) );
   IV110  g1379( .A(n5667), .Y(n6195) );
   IV110  g1380( .A(n5666), .Y(n5946) );
   IV110  g1381( .A(n5665), .Y(n5947) );
   BF003  g1382( .A1(n5789), .A2(n6561), .B1(n6181), .B2(
                           n6562), .Y(n6460) );
   BF003  g1383( .A1(n5788), .A2(n6459), .B1(n6083), .B2(
                           n6461), .Y(n6575) );
   EN210  g1384( .A(n6571), .B(n6550), .Y(n6576) );
   BF003  g1385( .A1(n5787), .A2(n6026), .B1(n6505), .B2(
                           n6027), .Y(n6103) );
   EN210  g1386( .A(n5413), .B(n6103), .Y(n5843) );
   EN210  g1387( .A(n5972), .B(n5971), .Y(n5970) );
   NA210  g1388( .A(A_2_port), .B(B_5_port), .Y(n5896) );
   NO210  g1389( .A(n6478), .B(n5234), .Y(n6330) );
   EX2B0  g1390( .A(n6125), .B(n5561), .Y(n5282) );
   NO210  g1391( .A(n6175), .B(n5232), .Y(n5899) );
   EN2B0  g1392( .A(n5987), .B(n5283), .Y(n5817) );
   NA210  g1393( .A(A_4_port), .B(B_4_port), .Y(n5640) );
   EX2B0  g1394( .A(n6426), .B(n5818), .Y(n5598) );
   NA210  g1395( .A(A_3_port), .B(B_5_port), .Y(n5641) );
   EN2B0  g1396( .A(n6435), .B(n5599), .Y(n6108) );
   BF003  g1397( .A1(n5254), .A2(n6465), .B1(n6078), .B2(
                           n5512), .Y(n6143) );
   BF003  g1398( .A1(n5253), .A2(n6556), .B1(n6079), .B2(
                           n5513), .Y(n6557) );
   EN210  g1399( .A(n6141), .B(n6557), .Y(n6144) );
   BF003  g1400( .A1(n5252), .A2(n5514), .B1(n6080), .B2(
                           n5515), .Y(n6553) );
   EN210  g1401( .A(n6142), .B(n6553), .Y(n6570) );
   BF003  g1402( .A1(n5251), .A2(n5516), .B1(n6081), .B2(
                           n5517), .Y(n5606) );
   IV110  g1403( .A(n5945), .Y(n5415) );
   EN210  g1404( .A(n6145), .B(n5606), .Y(n6573) );
   IV110  g1405( .A(n5942), .Y(n6369) );
   BF003  g1406( .A1(n5250), .A2(n5518), .B1(n6082), .B2(
                           n5520), .Y(n6572) );
   IV110  g1407( .A(n6564), .Y(n6563) );
   BF053  g1408( .A1(n6348), .A2(n6349), .B1(n5979), .B2(
                           n6044), .Y(n6562) );
   IV110  g1409( .A(n6562), .Y(n6561) );
   BF053  g1410( .A1(n6559), .A2(n6344), .B1(n5980), .B2(
                           n6042), .Y(n6560) );
   IV110  g1411( .A(n6560), .Y(n6135) );
   EX210  g1412( .A(n5943), .B(n6169), .Y(PRODUCT_27_port) );
   NA210  g1413( .A(B_0_port), .B(A_1_port), .Y(n6170) );
   NA210  g1414( .A(A_0_port), .B(B_1_port), .Y(n6171) );
   NO210  g1415( .A(n6170), .B(n6171), .Y(n5966) );
   AN210  g1416( .A(B_0_port), .B(A_2_port), .Y(n6243) );

endmodule

module rpl_add_n31_1

       ( A_30_port, A_29_port, A_28_port, A_27_port, A_26_port, A_25_port, 
         A_24_port, A_23_port, A_22_port, A_21_port, A_20_port, A_19_port, 
         A_18_port, A_17_port, A_16_port, A_15_port, A_14_port, A_13_port, 
         A_12_port, A_11_port, A_10_port, A_9_port, A_8_port, A_7_port, 
         A_6_port, A_5_port, A_4_port, A_3_port, A_2_port, A_1_port, A_0_port, 
         B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port, 
         B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port, 
         B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port, 
         B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port, 
         B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port, 
         SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
         SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
         SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
         SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
         SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, 
         SUM_6_port, SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port,
         SUM_0_port);

input A_30_port, A_29_port, A_28_port, A_27_port, A_26_port, A_25_port,
         A_24_port, A_23_port, A_22_port, A_21_port, A_20_port, A_19_port,
         A_18_port, A_17_port, A_16_port, A_15_port, A_14_port, A_13_port,
         A_12_port, A_11_port, A_10_port, A_9_port, A_8_port, A_7_port,
         A_6_port, A_5_port, A_4_port, A_3_port, A_2_port, A_1_port, A_0_port,
         B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port,
         B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port,
         B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port,
         B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
         B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port;

output   SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port,
         SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port,
         SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port,
         SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port,
         SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port,
         SUM_6_port, SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port,
         SUM_0_port;

   wire n188, n280, n189, n281, n282, n283, n284, n285, n286, n260, n287, 
      n261, n288, n262, n289, n263, n264, n265, n266, n240, n267, n241, n268, 
      n242, n269, n243, n244, n245, n246, n220, n247, n221, n248, n222, n249, 
      n223, n224, n225, n226, n200, n227, n201, n228, n202, n229, n203, n204, 
      n205, n206, n207, n208, n300, n209, n301, n302, n303, n304, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n290, n199, n291, n292, n293, 
      n294, n295, n296, n270, n297, n271, n298, n272, n299, n273, n274, n275, 
      n276, n250, n277, n251, n278, n252, n279, n253, n254, n255, n256, n230, 
      n257, n231, n258, n232, n259, n233, n234, n235, n236, n210, n237, n211, 
      n238, n212, n239, n213, n214, n215, n216, n217, n218, n219;

   BF003  g1( .A1(n302), .A2(n301), .B1(n216), .B2(n303), 
                           .Y(SUM_23_port) );
   BF003  g2( .A1(B_3_port), .A2(A_3_port), .B1(n217), .B2( 
                           n289), .Y(n198) );
   EX2B0  g3( .A(B_29_port), .B(A_29_port), .Y(n266) );
   BF003  g4( .A1(n253), .A2(n283), .B1(n256), .B2(n254), 
                           .Y(SUM_17_port) );
   BF003  g5( .A1(n298), .A2(n228), .B1(n300), .B2(n299), 
                           .Y(SUM_11_port) );
   IV110  g6( .A(n287), .Y(n238) );
   BF003  g7( .A1(n215), .A2(n200), .B1(A_2_port), .B2(
                           B_2_port), .Y(n291) );
   IV110  g8( .A(n286), .Y(n288) );
   BF003  g9( .A1(B_15_port), .A2(A_15_port), .B1(n281), .B2(
                           n237), .Y(n209) );
   BF003  g10( .A1(n286), .A2(n285), .B1(n288), .B2(n284), 
                           .Y(SUM_18_port) );
   BF003  g11( .A1(n274), .A2(n279), .B1(n278), .B2(n276), 
                           .Y(SUM_14_port) );
   BF003  g12( .A1(n251), .A2(n250), .B1(n211), .B2(n252), 
                           .Y(SUM_19_port) );
   BF003  g13( .A1(n289), .A2(n217), .B1(n291), .B2(n290), 
                           .Y(SUM_3_port) );
   IV110  g14( .A(n215), .Y(n248) );
   IV110  g15( .A(n193), .Y(n191) );
   EX2B0  g16( .A(B_10_port), .B(A_10_port), .Y(n226) );
   BF003  g17( .A1(n272), .A2(n271), .B1(n269), .B2(n273), 
                           .Y(SUM_28_port) );
   EX2B0  g18( .A(B_21_port), .B(A_21_port), .Y(n213) );
   BF003  g19( .A1(n200), .A2(n215), .B1(n249), .B2(n248), 
                           .Y(SUM_2_port) );
   BF003  g20( .A1(n208), .A2(n226), .B1(n255), .B2(n210), 
                           .Y(SUM_10_port) );
   BF003  g21( .A1(B_29_port), .A2(A_29_port), .B1(n266), .B2(
                           n235), .Y(n268) );
   IV110  g22( .A(n241), .Y(n237) );
   IV110  g23( .A(n283), .Y(n254) );
   EX2B0  g24( .A(B_9_port), .B(A_9_port), .Y(n225) );
   EX2B0  g25( .A(B_20_port), .B(A_20_port), .Y(n212) );
   BF003  g26( .A1(n204), .A2(n203), .B1(n218), .B2(n206), 
                           .Y(SUM_24_port) );
   IV110  g27( .A(n275), .Y(n201) );
   IV110  g28( .A(n217), .Y(n290) );
   IV110  g29( .A(n266), .Y(n260) );
   EX2B0  g30( .A(A_15_port), .B(B_15_port), .Y(n281) );
   EX2B0  g31( .A(B_26_port), .B(A_26_port), .Y(n265) );
   IV110  g32( .A(n255), .Y(n208) );
   IV110  g33( .A(n226), .Y(n210) );
   IV110  g34( .A(n214), .Y(n259) );
   IV110  g35( .A(n249), .Y(n200) );
   IV110  g36( .A(n281), .Y(n239) );
   EX2B0  g37( .A(A_14_port), .B(B_14_port), .Y(n279) );
   IV110  g38( .A(n216), .Y(n302) );
   BF003  g39( .A1(B_8_port), .A2(A_8_port), .B1(n224), .B2( 
                           n188), .Y(n232) );
   EX2B0  g40( .A(B_25_port), .B(A_25_port), .Y(n220) );
   IV110  g41( .A(n277), .Y(n246) );
   IV110  g42( .A(n262), .Y(n264) );
   IV110  g43( .A(n218), .Y(n204) );
   BF003  g44( .A1(B_26_port), .A2(A_26_port), .B1(n265), .B2(
                           n197), .Y(n242) );
   IV110  g45( .A(n228), .Y(n299) );
   BF003  g46( .A1(B_7_port), .A2(A_7_port), .B1(n223), .B2( 
                           n233), .Y(n190) );
   IV110  g47( .A(n220), .Y(n296) );
   BF003  g48( .A1(B_19_port), .A2(A_19_port), .B1(n211), .B2(
                           n252), .Y(n262) );
   IV110  g49( .A(n271), .Y(n273) );
   IV110  g50( .A(n280), .Y(n197) );
   IV110  g51( .A(n225), .Y(n231) );
   BF003  g52( .A1(B_6_port), .A2(A_6_port), .B1(n222), .B2( 
                           n191), .Y(n236) );
   BF003  g53( .A1(n296), .A2(n294), .B1(n220), .B2(n297), 
                           .Y(SUM_25_port) );
   IV110  g54( .A(n265), .Y(n195) );
   IV110  g55( .A(n250), .Y(n252) );
   BF003  g56( .A1(B_1_port), .A2(A_1_port), .B1(n293), .B2( 
                           A_0_port), .Y(n249) );
   BF003  g57( .A1(B_25_port), .A2(A_25_port), .B1(n220), .B2(
                           n297), .Y(n280) );
   BF003  g58( .A1(B_14_port), .A2(A_14_port), .B1(n279), .B2(
                           n274), .Y(n241) );
   BF003  g59( .A1(n284), .A2(n288), .B1(B_18_port), .B2(
                           A_18_port), .Y(n250) );
   BF003  g60( .A1(n245), .A2(n277), .B1(n247), .B2(n246), 
                           .Y(SUM_13_port) );
   NA210  g61( .A(B_0_port), .B(A_0_port), .Y(n292) );
   BF003  g62( .A1(B_13_port), .A2(A_13_port), .B1(n277), .B2(
                           n245), .Y(n278) );
   BF003  g63( .A1(n243), .A2(n242), .B1(n267), .B2(n244), 
                           .Y(SUM_27_port) );
   BF003  g64( .A1(n238), .A2(n221), .B1(n287), .B2(n240), 
                           .Y(SUM_5_port) );
   EX210  g65( .A(B_30_port), .B(A_30_port), .Y(n270) );
   IV110  g66( .A(n236), .Y(n233) );
   BF003  g67( .A1(B_12_port), .A2(A_12_port), .B1(n275), .B2(
                           n199), .Y(n247) );
   EX2B0  g68( .A(B_28_port), .B(A_28_port), .Y(n269) );
   IV110  g69( .A(n257), .Y(n261) );
   BF003  g70( .A1(n194), .A2(n219), .B1(n198), .B2(n196), 
                           .Y(SUM_4_port) );
   BF003  g71( .A1(n233), .A2(n223), .B1(n236), .B2(n234), 
                           .Y(SUM_7_port) );
   IV110  g72( .A(n190), .Y(n188) );
   EX2B0  g73( .A(B_27_port), .B(A_27_port), .Y(n267) );
   BF003  g74( .A1(n237), .A2(n281), .B1(n241), .B2(n239), 
                           .Y(SUM_15_port) );
   BF003  g75( .A1(n191), .A2(n222), .B1(n193), .B2(n192), 
                           .Y(SUM_6_port) );
   IV110  g76( .A(n291), .Y(n289) );
   BF003  g77( .A1(n230), .A2(n225), .B1(n232), .B2(n231), 
                           .Y(SUM_9_port) );
   IV110  g78( .A(n209), .Y(n205) );
   BF003  g80( .A1(B_5_port), .A2(A_5_port), .B1(n221), .B2( 
                           n238), .Y(n193) );
   EX2B0  g81( .A(A_19_port), .B(B_19_port), .Y(n211) );
   BF003  g82( .A1(n199), .A2(n275), .B1(n202), .B2(n201), 
                           .Y(SUM_12_port) );
   BF003  g83( .A1(n260), .A2(n258), .B1(n266), .B2(n235), 
                           .Y(SUM_29_port) );
   IV110  g84( .A(n198), .Y(n194) );
   EX2B0  g85( .A(B_23_port), .B(A_23_port), .Y(n216) );
   IV110  g86( .A(n256), .Y(n253) );
   BF003  g87( .A1(n263), .A2(n262), .B1(n212), .B2(n264), 
                           .Y(SUM_20_port) );
   BF003  g88( .A1(n205), .A2(n282), .B1(n209), .B2(n207), 
                           .Y(SUM_16_port) );
   BF003  g89( .A1(B_28_port), .A2(A_28_port), .B1(n269), .B2(
                           n273), .Y(n258) );
   BF003  g90( .A1(n195), .A2(n280), .B1(n265), .B2(n197), 
                           .Y(SUM_26_port) );
   IV110  g91( .A(n247), .Y(n245) );
   IV110  g92( .A(n219), .Y(n196) );
   EX2B0  g93( .A(A_11_port), .B(B_11_port), .Y(n228) );
   EX2B0  g94( .A(B_22_port), .B(A_22_port), .Y(n214) );
   BF003  g95( .A1(n259), .A2(n257), .B1(n214), .B2(n261), 
                           .Y(SUM_22_port) );
   IV110  g96( .A(n258), .Y(n235) );
   IV110  g97( .A(n278), .Y(n274) );
   IV110  g98( .A(n300), .Y(n298) );
   IV110  g99( .A(n224), .Y(n189) );
   IV110  g100( .A(n284), .Y(n285) );
   EX2B0  g101( .A(A_13_port), .B(B_13_port), .Y(n277) );
   EX2B0  g102( .A(B_24_port), .B(A_24_port), .Y(n218) );
   BF003  g103( .A1(B_27_port), .A2(A_27_port), .B1(n267), .B2(
                           n244), .Y(n271) );
   IV110  g104( .A(n202), .Y(n199) );
   EX2B0  g105( .A(B_18_port), .B(A_18_port), .Y(n284) );
   IV110  g106( .A(n222), .Y(n192) );
   IV110  g107( .A(n282), .Y(n207) );
   IV110  g108( .A(n211), .Y(n251) );
   IV110  g109( .A(n223), .Y(n234) );
   IV110  g110( .A(n294), .Y(n297) );
   EX2B0  g111( .A(A_12_port), .B(B_12_port), .Y(n275) );
   IV110  g112( .A(n267), .Y(n243) );
   BF003  g113( .A1(B_17_port), .A2(A_17_port), .B1(n283), .B2(
                           n253), .Y(n286) );
   EX2B0  g114( .A(B_17_port), .B(A_17_port), .Y(n283) );
   BF003  g115( .A1(B_24_port), .A2(A_24_port), .B1(n218), .B2(
                           n206), .Y(n294) );
   IV110  g116( .A(n279), .Y(n276) );
   BF003  g117( .A1(B_16_port), .A2(A_16_port), .B1(n282), .B2(
                           n205), .Y(n256) );
   IV110  g118( .A(n221), .Y(n240) );
   IV110  g119( .A(n203), .Y(n206) );
   IV110  g120( .A(n269), .Y(n272) );
   BF003  g121( .A1(B_23_port), .A2(A_23_port), .B1(n216), .B2(
                           n303), .Y(n203) );
   EX2B0  g122( .A(A_16_port), .B(B_16_port), .Y(n282) );
   IV110  g123( .A(n301), .Y(n303) );
   AN210  g124( .A(n295), .B(B_0_port), .Y(n293) );
   IV110  g125( .A(n232), .Y(n230) );
   EX2B0  g126( .A(B_5_port), .B(A_5_port), .Y(n221) );
   BF003  g127( .A1(B_22_port), .A2(A_22_port), .B1(n214), .B2(
                           n261), .Y(n301) );
   BF003  g128( .A1(B_11_port), .A2(A_11_port), .B1(n228), .B2(
                           n298), .Y(n202) );
   EX2B0  g129( .A(A_4_port), .B(B_4_port), .Y(n219) );
   EX2B0  g130( .A(B_8_port), .B(A_8_port), .Y(n224) );
   BF003  g131( .A1(B_21_port), .A2(A_21_port), .B1(n213), .B2(
                           n229), .Y(n257) );
   EX2B0  g132( .A(A_3_port), .B(B_3_port), .Y(n217) );
   EX2B0  g133( .A(B_7_port), .B(A_7_port), .Y(n223) );
   EX210  g134( .A(B_0_port), .B(A_0_port), .Y(SUM_0_port) );
   EX2B0  g135( .A(A_2_port), .B(B_2_port), .Y(n215) );
   BF003  g136( .A1(B_10_port), .A2(A_10_port), .B1(n226), .B2(
                           n208), .Y(n300) );
   EX2B0  g137( .A(A_1_port), .B(B_1_port), .Y(n295) );
   EX2B0  g138( .A(A_6_port), .B(B_6_port), .Y(n222) );
   IV110  g139( .A(n304), .Y(n229) );
   IV110  g140( .A(n212), .Y(n263) );
   EN210  g141( .A(n295), .B(n292), .Y(SUM_1_port) );
   BF003  g142( .A1(n188), .A2(n224), .B1(n190), .B2(n189), 
                           .Y(SUM_8_port) );
   IV110  g143( .A(n213), .Y(n227) );
   BF003  g144( .A1(B_9_port), .A2(A_9_port), .B1(n225), .B2( 
                           n230), .Y(n255) );
   BF003  g145( .A1(n227), .A2(n304), .B1(n213), .B2(n229), 
                           .Y(SUM_21_port) );
   BF003  g146( .A1(B_20_port), .A2(A_20_port), .B1(n212), .B2(
                           n264), .Y(n304) );
   BF003  g147( .A1(B_4_port), .A2(A_4_port), .B1(n219), .B2( 
                           n194), .Y(n287) );
   IV110  g148( .A(n242), .Y(n244) );
   EN210  g149( .A(n270), .B(n268), .Y(SUM_30_port) );

endmodule

module multx16 

       ( a_15_port, a_14_port, a_13_port, a_12_port, a_11_port, a_10_port, 
         a_9_port, a_8_port, a_7_port, a_6_port, a_5_port, a_4_port, a_3_port, 
         a_2_port, a_1_port, a_0_port, b_15_port, b_14_port, b_13_port, 
         b_12_port, b_11_port, b_10_port, b_9_port, b_8_port, b_7_port, 
         b_6_port, b_5_port, b_4_port, b_3_port, b_2_port, b_1_port, b_0_port, 
         c_15_port, c_14_port, c_13_port, c_12_port, c_11_port, c_10_port, 
         c_9_port, c_8_port, c_7_port, c_6_port, c_5_port, c_4_port, c_3_port, 
         c_2_port, c_1_port, c_0_port, d_15_port, d_14_port, d_13_port, 
         d_12_port, d_11_port, d_10_port, d_9_port, d_8_port, d_7_port, 
         d_6_port, d_5_port, d_4_port, d_3_port, d_2_port, d_1_port, d_0_port, 
         sel_3_port, sel_2_port, sel_1_port, sel_0_port,  
         y_30_port, y_29_port, y_28_port, y_27_port, y_26_port, y_25_port, 
         y_24_port, y_23_port, y_22_port, y_21_port, y_20_port, y_19_port, 
         y_18_port, y_17_port, y_16_port, y_15_port, y_14_port, y_13_port, 
         y_12_port, y_11_port, y_10_port, y_9_port, y_8_port, y_7_port, 
         y_6_port, y_5_port, y_4_port, y_3_port, y_2_port, y_1_port, y_0_port );

input a_15_port, a_14_port, a_13_port, a_12_port, a_11_port, a_10_port,
         a_9_port, a_8_port, a_7_port, a_6_port, a_5_port, a_4_port, a_3_port,
         a_2_port, a_1_port, a_0_port, b_15_port, b_14_port, b_13_port,
         b_12_port, b_11_port, b_10_port, b_9_port, b_8_port, b_7_port,
         b_6_port, b_5_port, b_4_port, b_3_port, b_2_port, b_1_port, b_0_port,
         c_15_port, c_14_port, c_13_port, c_12_port, c_11_port, c_10_port,
         c_9_port, c_8_port, c_7_port, c_6_port, c_5_port, c_4_port, c_3_port,
         c_2_port, c_1_port, c_0_port, d_15_port, d_14_port, d_13_port,
         d_12_port, d_11_port, d_10_port, d_9_port, d_8_port, d_7_port,
         d_6_port, d_5_port, d_4_port, d_3_port, d_2_port, d_1_port, d_0_port,
         sel_3_port, sel_2_port, sel_1_port, sel_0_port;

output y_30_port, y_29_port, y_28_port, y_27_port, y_26_port, y_25_port,
         y_24_port, y_23_port, y_22_port, y_21_port, y_20_port, y_19_port,
         y_18_port, y_17_port, y_16_port, y_15_port, y_14_port, y_13_port,
         y_12_port, y_11_port, y_10_port, y_9_port, y_8_port, y_7_port,
         y_6_port, y_5_port, y_4_port, y_3_port, y_2_port, y_1_port, y_0_port;
 

   wire y2_5_port, y2_7_port, y2_9_port, n25, n26, y1_8_port, y1_6_port, 
      y1_4_port, y2_21_port, y1_21_port, y1_2_port, y2_23_port, y1_23_port, 
      Logic0, y1_0_port, y2_11_port, y1_11_port, y2_25_port, y1_25_port, 
      y2_13_port, y1_13_port, y2_27_port, y1_27_port, y2_15_port, y1_15_port, 
      y2_29_port, y1_29_port, y2_17_port, y1_17_port, y2_19_port, y1_19_port, 
      y2_0_port, y2_2_port, y2_4_port, y2_6_port, y2_8_port, y1_9_port, 
      y1_7_port, y2_30_port, y1_30_port, y1_5_port, y2_20_port, y1_20_port, 
      y1_3_port, y2_22_port, y1_22_port, y1_1_port, y2_10_port, y1_10_port, 
      y2_24_port, y1_24_port, y2_12_port, y1_12_port, y2_26_port, y1_26_port, 
      y2_14_port, y1_14_port, y2_28_port, y1_28_port, y2_16_port, y1_16_port, 
      y2_18_port, y1_18_port, y2_1_port, y2_3_port;

   rpl_add_n31_1   m1  	 ( .A_30_port(y2_30_port), .A_29_port( 
                           y2_29_port), .A_28_port(y2_28_port), .A_27_port(
                           y2_27_port), .A_26_port(y2_26_port), .A_25_port(
                           y2_25_port), .A_24_port(y2_24_port), .A_23_port(
                           y2_23_port), .A_22_port(y2_22_port), .A_21_port(
                           y2_21_port), .A_20_port(y2_20_port), .A_19_port(
                           y2_19_port), .A_18_port(y2_18_port), .A_17_port(
                           y2_17_port), .A_16_port(y2_16_port), .A_15_port(
                           y2_15_port), .A_14_port(y2_14_port), .A_13_port(
                           y2_13_port), .A_12_port(y2_12_port), .A_11_port(
                           y2_11_port), .A_10_port(y2_10_port), .A_9_port(
                           y2_9_port), .A_8_port(y2_8_port), .A_7_port(
                           y2_7_port), .A_6_port(y2_6_port), .A_5_port(
                           y2_5_port), .A_4_port(y2_4_port), .A_3_port(
                           y2_3_port), .A_2_port(y2_2_port), .A_1_port(
                           y2_1_port), .A_0_port(y2_0_port), .B_30_port(
                           y1_30_port), .B_29_port(y1_29_port), .B_28_port(
                           y1_28_port), .B_27_port(y1_27_port), .B_26_port(
                           y1_26_port), .B_25_port(y1_25_port), .B_24_port(
                           y1_24_port), .B_23_port(y1_23_port), .B_22_port(
                           y1_22_port), .B_21_port(y1_21_port), .B_20_port(
                           y1_20_port), .B_19_port(y1_19_port), .B_18_port(
                           y1_18_port), .B_17_port(y1_17_port), .B_16_port(
                           y1_16_port), .B_15_port(y1_15_port), .B_14_port(
                           y1_14_port), .B_13_port(y1_13_port), .B_12_port(
                           y1_12_port), .B_11_port(y1_11_port), .B_10_port(
                           y1_10_port), .B_9_port(y1_9_port), .B_8_port(
                           y1_8_port), .B_7_port(y1_7_port), .B_6_port(
                           y1_6_port), .B_5_port(y1_5_port), .B_4_port(
                           y1_4_port), .B_3_port(y1_3_port), .B_2_port(
                           y1_2_port), .B_1_port(y1_1_port), .B_0_port(
                           y1_0_port), .SUM_30_port(y_30_port), .SUM_29_port(
                           y_29_port), .SUM_28_port(y_28_port), .SUM_27_port(
                           y_27_port), .SUM_26_port(y_26_port), .SUM_25_port(
                           y_25_port), .SUM_24_port(y_24_port), .SUM_23_port(
                           y_23_port), .SUM_22_port(y_22_port), .SUM_21_port(
                           y_21_port), .SUM_20_port(y_20_port), .SUM_19_port(
                           y_19_port), .SUM_18_port(y_18_port), .SUM_17_port(
                           y_17_port), .SUM_16_port(y_16_port), .SUM_15_port(
                           y_15_port), .SUM_14_port(y_14_port), .SUM_13_port(
                           y_13_port), .SUM_12_port(y_12_port), .SUM_11_port(
                           y_11_port), .SUM_10_port(y_10_port), .SUM_9_port(
                           y_9_port), .SUM_8_port(y_8_port), .SUM_7_port(
                           y_7_port), .SUM_6_port(y_6_port), .SUM_5_port(
                           y_5_port), .SUM_4_port(y_4_port), .SUM_3_port(
                           y_3_port), .SUM_2_port(y_2_port), .SUM_1_port(
                           y_1_port), .SUM_0_port(y_0_port));

   csa_mult_n17_m17_1  m2 ( .A_16_port(Logic0), .A_15_port(
                           b_15_port), .A_14_port(b_14_port), .A_13_port(
                           b_13_port), .A_12_port(b_12_port), .A_11_port(
                           b_11_port), .A_10_port(b_10_port), .A_9_port(
                           b_9_port), .A_8_port(b_8_port), .A_7_port(b_7_port
                           ), .A_6_port(b_6_port), .A_5_port(b_5_port), 
                           .A_4_port(b_4_port), .A_3_port(b_3_port), .A_2_port
                          (b_2_port), .A_1_port(b_1_port), .A_0_port(
                           b_0_port), .B_16_port(Logic0), .B_15_port(
                           a_15_port), .B_14_port(a_14_port), .B_13_port(
                           a_13_port), .B_12_port(a_12_port), .B_11_port(
                           a_11_port), .B_10_port(a_10_port), .B_9_port(
                           a_9_port), .B_8_port(a_8_port), .B_7_port(a_7_port
                           ), .B_6_port(a_6_port), .B_5_port(a_5_port), 
                           .B_4_port(a_4_port), .B_3_port(a_3_port), .B_2_port
                          (a_2_port), .B_1_port(a_1_port), .B_0_port(
                           a_0_port), .CTL(n25), .PRODUCT_33_port(open), 
                           .PRODUCT_32_port(open), .PRODUCT_31_port(open), 
                           .PRODUCT_30_port(y1_30_port), .PRODUCT_29_port(
                           y1_29_port), .PRODUCT_28_port(y1_28_port), 
                           .PRODUCT_27_port(y1_27_port), .PRODUCT_26_port(
                           y1_26_port), .PRODUCT_25_port(y1_25_port), 
                           .PRODUCT_24_port(y1_24_port), .PRODUCT_23_port(
                           y1_23_port), .PRODUCT_22_port(y1_22_port), 
                           .PRODUCT_21_port(y1_21_port), .PRODUCT_20_port(
                           y1_20_port), .PRODUCT_19_port(y1_19_port), 
                           .PRODUCT_18_port(y1_18_port), .PRODUCT_17_port(
                           y1_17_port), .PRODUCT_16_port(y1_16_port), 
                           .PRODUCT_15_port(y1_15_port), .PRODUCT_14_port(
                           y1_14_port), .PRODUCT_13_port(y1_13_port), 
                           .PRODUCT_12_port(y1_12_port), .PRODUCT_11_port(
                           y1_11_port), .PRODUCT_10_port(y1_10_port), 
                           .PRODUCT_9_port(y1_9_port), .PRODUCT_8_port(
                           y1_8_port), .PRODUCT_7_port(y1_7_port), 
                           .PRODUCT_6_port(y1_6_port), .PRODUCT_5_port(
                           y1_5_port), .PRODUCT_4_port(y1_4_port), 
                           .PRODUCT_3_port(y1_3_port), .PRODUCT_2_port(
                           y1_2_port), .PRODUCT_1_port(y1_1_port), 
                           .PRODUCT_0_port(y1_0_port));

   csa_mult_n17_m17_2  m3 ( .A_16_port(Logic0), .A_15_port(
                           d_15_port), .A_14_port(d_14_port), .A_13_port(
                           d_13_port), .A_12_port(d_12_port), .A_11_port(
                           d_11_port), .A_10_port(d_10_port), .A_9_port(
                           d_9_port), .A_8_port(d_8_port), .A_7_port(d_7_port
                           ), .A_6_port(d_6_port), .A_5_port(d_5_port), 
                           .A_4_port(d_4_port), .A_3_port(d_3_port), .A_2_port
                          (d_2_port), .A_1_port(d_1_port), .A_0_port(
                           d_0_port), .B_16_port(Logic0), .B_15_port(
                           c_15_port), .B_14_port(c_14_port), .B_13_port(
                           c_13_port), .B_12_port(c_12_port), .B_11_port(
                           c_11_port), .B_10_port(c_10_port), .B_9_port(
                           c_9_port), .B_8_port(c_8_port), .B_7_port(c_7_port
                           ), .B_6_port(c_6_port), .B_5_port(c_5_port), 
                           .B_4_port(c_4_port), .B_3_port(c_3_port), .B_2_port
                          (c_2_port), .B_1_port(c_1_port), .B_0_port(
                           c_0_port), .CTL(n26), .PRODUCT_33_port(open), 
                           .PRODUCT_32_port(open), .PRODUCT_31_port(open), 
                           .PRODUCT_30_port(y2_30_port), .PRODUCT_29_port(
                           y2_29_port), .PRODUCT_28_port(y2_28_port), 
                           .PRODUCT_27_port(y2_27_port), .PRODUCT_26_port(
                           y2_26_port), .PRODUCT_25_port(y2_25_port), 
                           .PRODUCT_24_port(y2_24_port), .PRODUCT_23_port(
                           y2_23_port), .PRODUCT_22_port(y2_22_port), 
                           .PRODUCT_21_port(y2_21_port), .PRODUCT_20_port(
                           y2_20_port), .PRODUCT_19_port(y2_19_port), 
                           .PRODUCT_18_port(y2_18_port), .PRODUCT_17_port(
                           y2_17_port), .PRODUCT_16_port(y2_16_port), 
                           .PRODUCT_15_port(y2_15_port), .PRODUCT_14_port(
                           y2_14_port), .PRODUCT_13_port(y2_13_port), 
                           .PRODUCT_12_port(y2_12_port), .PRODUCT_11_port(
                           y2_11_port), .PRODUCT_10_port(y2_10_port), 
                           .PRODUCT_9_port(y2_9_port), .PRODUCT_8_port(
                           y2_8_port), .PRODUCT_7_port(y2_7_port), 
                           .PRODUCT_6_port(y2_6_port), .PRODUCT_5_port(
                           y2_5_port), .PRODUCT_4_port(y2_4_port), 
                           .PRODUCT_3_port(y2_3_port), .PRODUCT_2_port(
                           y2_2_port), .PRODUCT_1_port(y2_1_port), 
                           .PRODUCT_0_port(y2_0_port));
TO010  m4 ( .HI(open), .LO(Logic0));
TO010  m5 ( .HI(n25), .LO(open));
TO010  m6 ( .HI(n26), .LO(open));
and	test1 ( testout, sel_0_port, sel_1_port, sel_2_port, sel_3_port);


endmodule

// End of public domain circuit
