module zero ( LO );

// Verilog Port Declaration section

   output LO;


// Verilog Structure section (in terms of gate prims)


           buf  #1 ( LO , 1'b0 ) ;

endmodule
